magic
tech sky130B
magscale 1 2
timestamp 1713529395
<< error_p >>
rect 566 7884 572 7896
rect 804 7884 810 7896
rect 578 7872 590 7878
rect 786 7872 798 7878
<< error_s >>
rect 23816 11208 23822 11210
rect 23893 11208 23899 11210
rect 23816 11205 23830 11208
rect 23885 11205 23899 11208
rect 23816 11204 23822 11205
rect 23893 11204 23899 11205
rect 23810 11199 23905 11204
rect 23810 11198 23821 11199
rect 23674 11053 23730 11197
rect 23812 11190 23821 11198
rect 23894 11198 23905 11199
rect 23894 11190 23903 11198
rect 23816 11135 23821 11190
rect 23812 11127 23821 11135
rect 23810 11126 23821 11127
rect 23894 11127 23903 11135
rect 23894 11126 23905 11127
rect 23810 11121 23905 11126
rect 23816 11120 23822 11121
rect 23893 11120 23899 11121
rect 23816 11117 23830 11120
rect 23885 11117 23899 11120
rect 23816 11115 23822 11117
rect 23893 11115 23899 11117
rect 23674 11003 24018 11053
rect 23674 10979 23730 11003
rect 23638 10943 24078 10973
rect 23354 10659 23730 10877
rect 27542 10766 27548 10778
rect 27624 10766 27630 10778
rect 27554 10754 27566 10760
rect 27606 10754 27618 10760
rect 27606 10188 27618 10194
rect 27624 10170 27630 10182
rect 27624 10118 27630 10130
rect 27606 10106 27618 10112
rect 27970 9616 27982 9622
rect 27958 9598 27964 9610
rect 26999 9376 27074 9379
rect 28226 9376 28289 9379
rect 26999 9342 27108 9345
rect 28192 9342 28289 9345
rect 28400 8510 28412 8516
rect 28418 8492 28424 8504
rect 28418 8284 28424 8296
rect 41656 8282 41662 8294
rect 41894 8282 41900 8294
rect 28400 8272 28412 8278
rect 41668 8270 41680 8276
rect 41876 8270 41888 8276
rect 47593 8240 47599 8252
rect 47697 8240 47703 8252
rect 47605 8228 47617 8234
rect 47679 8228 47691 8234
rect 46966 8157 46978 8163
rect 46954 8139 46960 8151
rect 46954 8087 46960 8099
rect 46966 8075 46978 8081
rect 10360 7992 10372 7998
rect 10348 7974 10354 7986
rect 10348 7922 10354 7934
rect 10360 7910 10372 7916
rect 6503 7842 6509 7854
rect 6607 7842 6613 7854
rect 6515 7830 6527 7836
rect 6589 7830 6601 7836
rect 5876 7759 5888 7765
rect 5864 7741 5870 7753
rect 12344 7704 12356 7710
rect 12396 7704 12408 7710
rect 5864 7689 5870 7701
rect 12332 7686 12338 7698
rect 12414 7686 12420 7698
rect 5876 7677 5888 7683
rect 19950 7378 19962 7384
rect 19938 7360 19944 7372
rect 19938 7308 19944 7320
rect 19950 7296 19962 7302
rect 47590 6380 47608 6386
rect 47670 6380 47688 6386
rect 47584 6362 47590 6380
rect 47688 6362 47694 6380
rect 47584 6282 47590 6300
rect 47688 6282 47694 6300
rect 47590 6276 47608 6282
rect 47670 6276 47688 6282
rect 34286 6096 34292 6102
rect 34512 6096 34518 6102
rect 46538 6096 46544 6108
rect 46620 6096 46626 6108
rect 48960 6098 48978 6104
rect 49018 6098 49036 6104
rect 34280 6090 34286 6096
rect 34518 6090 34524 6096
rect 46550 6084 46562 6090
rect 46602 6084 46614 6090
rect 48954 6080 48960 6098
rect 49036 6080 49042 6098
rect 48954 6022 48960 6040
rect 49036 6022 49042 6040
rect 48960 6016 48978 6022
rect 49018 6016 49036 6022
rect 6500 5982 6518 5988
rect 6580 5982 6598 5988
rect 6494 5964 6500 5982
rect 6598 5964 6604 5982
rect 6494 5884 6500 5902
rect 6598 5884 6604 5902
rect 6500 5878 6518 5884
rect 6580 5878 6598 5884
rect 12753 5864 12756 5870
rect 34280 5864 34286 5870
rect 34518 5864 34524 5870
rect 34286 5858 34292 5864
rect 34512 5858 34518 5864
rect 12765 5846 12768 5858
rect 5448 5698 5454 5710
rect 5530 5698 5536 5710
rect 7876 5700 7888 5706
rect 5460 5686 5472 5692
rect 5512 5686 5524 5692
rect 7864 5682 7870 5694
rect 7864 5630 7870 5642
rect 12765 5638 12768 5650
rect 12744 5626 12756 5632
rect 7876 5618 7888 5624
rect 9756 5387 9757 5393
rect 9744 5369 9750 5381
rect 9756 5320 9818 5346
rect 9718 5282 9730 5308
rect 9796 5282 9830 5308
rect 9696 4774 9730 4784
rect 9796 4774 9818 4784
rect 9717 4736 9780 4746
rect 9705 4687 9711 4699
rect 9786 4687 9792 4699
rect 9717 4675 9719 4681
rect 9778 4675 9780 4681
rect 47338 4525 47344 4537
rect 47420 4525 47426 4537
rect 47350 4513 47362 4519
rect 47402 4513 47414 4519
rect 6248 4127 6254 4139
rect 6330 4127 6336 4139
rect 6260 4115 6272 4121
rect 6312 4115 6324 4121
rect 9719 4020 9778 4021
rect 9696 3986 9778 4020
rect 9796 3986 9816 4020
rect 9719 3962 9778 3986
rect 47338 3053 47344 3065
rect 47420 3053 47426 3065
rect 47350 3041 47362 3047
rect 47402 3041 47414 3047
rect 9719 2732 9778 2735
rect 9696 2698 9778 2732
rect 9796 2698 9816 2732
rect 9719 2676 9778 2698
rect 6248 2655 6254 2667
rect 6330 2655 6336 2667
rect 6260 2643 6272 2649
rect 6312 2643 6324 2649
rect 46794 2284 46806 2290
rect 46812 2266 46818 2278
rect 46812 2214 46818 2226
rect 46794 2202 46806 2208
rect 5704 1886 5716 1892
rect 5722 1868 5728 1880
rect 5722 1816 5728 1828
rect 5704 1804 5716 1810
rect 9719 1449 9778 1474
rect 9696 1415 9778 1449
rect 9696 1410 9730 1415
rect 9796 1410 9816 1444
rect 11322 1280 11530 1488
rect 11907 1296 11923 1307
rect 13201 1296 13211 1315
rect 14486 1296 14499 1315
rect 15776 1296 15787 1315
rect 17062 1296 17075 1315
rect 18354 1296 18363 1315
rect 19642 1296 19651 1315
rect 20927 1296 20939 1315
rect 13286 1288 13298 1289
rect 21012 1283 21024 1289
rect 11907 1196 11923 1230
rect 11945 1222 11961 1269
rect 13201 1196 13211 1230
rect 13239 1214 13249 1277
rect 13304 1276 13310 1277
rect 14486 1196 14499 1230
rect 14524 1217 14537 1277
rect 15776 1196 15787 1230
rect 15814 1218 15825 1277
rect 17062 1196 17075 1230
rect 17100 1218 17113 1277
rect 18354 1196 18363 1230
rect 18392 1218 18401 1277
rect 19642 1196 19651 1230
rect 19680 1218 19689 1277
rect 20927 1196 20939 1230
rect 20965 1218 20977 1277
rect 21030 1265 21036 1277
rect 21030 1218 21036 1230
rect 21012 1206 21024 1212
rect 26432 -2344 26451 -1987
rect 26384 -2345 26393 -2344
rect 26431 -2345 26451 -2344
rect 26382 -2348 26400 -2345
rect 26424 -2348 26451 -2345
rect 26379 -2349 26445 -2348
rect 26374 -2351 26380 -2349
rect 26382 -2351 26400 -2349
rect 26424 -2351 26442 -2349
rect 26374 -2369 26382 -2351
rect 26442 -2353 26448 -2351
rect 26442 -2362 26449 -2353
rect 26442 -2369 26448 -2362
rect 26374 -2393 26380 -2369
rect 26374 -2411 26382 -2393
rect 26442 -2400 26448 -2393
rect 26442 -2409 26449 -2400
rect 26442 -2411 26448 -2409
rect 26374 -2413 26380 -2411
rect 26382 -2413 26400 -2411
rect 26424 -2413 26442 -2411
rect 26379 -2414 26445 -2413
rect 26382 -2417 26400 -2414
rect 26424 -2417 26442 -2414
rect 26384 -2418 26393 -2417
rect 26431 -2418 26440 -2417
<< locali >>
rect 27970 10694 28100 10758
rect 26913 9345 26999 9462
rect 28289 9345 28375 9487
rect 26913 9259 28375 9345
rect 8944 8066 11011 8152
rect 11097 8066 13146 8152
rect 19192 7740 19905 7826
rect 20009 7740 20922 7826
rect 10178 4131 10250 4625
rect 10347 4267 10414 4524
rect 10179 2867 10251 3072
rect 10345 2973 10412 3236
rect 10179 1579 10251 1782
rect 10347 1741 10414 1927
rect 9726 300 9782 582
rect 10717 300 10828 2328
rect 13497 1722 13513 1809
rect 13661 1722 13678 1809
rect 12072 1579 12304 1651
rect 13360 1579 13577 1651
rect 14648 1579 14867 1651
rect 15936 1579 16159 1651
rect 17224 1578 17432 1650
rect 18512 1578 18731 1650
rect 19800 1579 20009 1651
rect 21088 1579 21289 1651
rect 12249 300 12365 642
rect 13534 300 13650 642
rect 14833 300 14949 642
rect 16117 300 16233 642
rect 17402 300 17518 642
rect 18687 300 18803 642
rect 19976 300 20092 642
rect 26913 311 26999 9259
rect 35042 5592 38198 5812
rect 28192 311 28412 1236
rect 26805 310 32886 311
rect 36278 310 36498 5592
rect 45593 310 45895 707
rect 8100 9 21424 300
rect 8103 0 21424 9
rect 21124 -2297 21424 0
rect 26805 8 45895 310
rect 26805 -2297 27108 8
rect 21124 -2334 26204 -2297
rect 26504 -2334 27108 -2297
rect 21124 -2357 27108 -2334
rect 21124 -2405 26388 -2357
rect 26436 -2405 27108 -2357
rect 21124 -2597 27108 -2405
rect 26805 -2598 27108 -2597
<< viali >>
rect 27554 10766 27618 10830
rect 26998 10124 27050 10176
rect 27554 10118 27618 10182
rect 27970 9546 28034 9610
rect 11011 8066 11097 8152
rect 10360 7922 10424 7986
rect 12756 7922 12820 7986
rect 19905 7722 20009 7826
rect 9763 7650 9812 7699
rect 12344 7634 12408 7698
rect 20558 7461 20610 7513
rect 19950 7308 20014 7372
rect 5894 5620 5946 5672
rect 7876 5630 7940 5694
rect 11316 5638 11536 5858
rect 12533 5638 12756 5858
rect 9756 5320 9818 5381
rect 9717 4687 9780 4746
rect 9719 3962 9778 4021
rect 9719 2676 9778 2735
rect 9719 1415 9778 1474
rect 11322 1280 11530 1488
rect 11945 1222 11992 1269
rect 13239 1214 13298 1277
rect 14524 1217 14584 1277
rect 15814 1218 15873 1277
rect 17100 1218 17159 1277
rect 18392 1218 18451 1277
rect 19680 1218 19739 1277
rect 20965 1218 21024 1277
rect 28192 8284 28412 8504
rect 33159 5877 33370 6088
rect 34292 5870 34512 6090
rect 46971 6018 47020 6067
rect 48966 6028 49030 6092
rect 39156 5597 39359 5800
rect 26388 -2405 26436 -2357
<< metal1 >>
rect 20904 11858 29116 12158
rect 20904 8700 21204 11858
rect 23400 11490 27618 11500
rect 23400 11436 27554 11490
rect 23400 11199 23464 11436
rect 27548 11426 27554 11436
rect 27618 11426 27624 11490
rect 7800 8400 21204 8700
rect 21623 11126 23821 11199
rect 23894 11126 23900 11199
rect 11011 8158 11097 8400
rect 10999 8152 11109 8158
rect 10999 8066 11011 8152
rect 11097 8066 11109 8152
rect 10999 8060 11109 8066
rect 10354 7986 10430 7992
rect 12750 7987 12826 7992
rect 11045 7986 11109 7987
rect 12750 7986 13916 7987
rect 10354 7922 10360 7986
rect 10424 7922 12756 7986
rect 12820 7922 13916 7986
rect 10354 7916 10430 7922
rect 9757 7699 9818 7711
rect 9757 7650 9763 7699
rect 9812 7650 9818 7699
rect 9568 6879 9632 6885
rect 7460 6224 9370 6288
rect 9434 6224 9440 6288
rect 7244 6100 7308 6106
rect 9568 6100 9632 6815
rect 5888 6036 7244 6100
rect 7694 6036 7700 6100
rect 7764 6036 9632 6100
rect 5888 5672 5952 6036
rect 7244 6030 7308 6036
rect 9757 5866 9818 7650
rect 11045 7056 11109 7922
rect 12750 7921 13916 7922
rect 12750 7916 12826 7921
rect 12338 7698 12414 7704
rect 12338 7634 12344 7698
rect 12408 7634 12414 7698
rect 13850 7686 13916 7921
rect 19905 7832 20009 8400
rect 19893 7826 20021 7832
rect 19893 7722 19905 7826
rect 20009 7722 20021 7826
rect 19893 7716 20021 7722
rect 12338 7628 12414 7634
rect 10548 6988 10554 7056
rect 10618 6992 11109 7056
rect 10618 6988 10624 6992
rect 9980 6879 10044 6885
rect 12344 6879 12408 7628
rect 13838 7622 18950 7686
rect 13850 7619 13916 7622
rect 18886 7519 18950 7622
rect 20552 7519 20616 7525
rect 18886 7513 20616 7519
rect 18886 7461 20558 7513
rect 20610 7461 20616 7513
rect 18886 7455 20616 7461
rect 20552 7449 20616 7455
rect 21623 7417 21696 11126
rect 27554 10836 27618 11426
rect 27548 10830 27624 10836
rect 27548 10766 27554 10830
rect 27618 10766 27624 10830
rect 27548 10760 27624 10766
rect 27548 10182 27624 10188
rect 26986 10176 27554 10182
rect 26986 10124 26998 10176
rect 27050 10124 27554 10176
rect 26986 10118 27554 10124
rect 27618 10118 27624 10182
rect 27548 10112 27624 10118
rect 28816 9744 29116 11858
rect 28816 9708 45822 9744
rect 27964 9614 28040 9616
rect 27964 9610 28186 9614
rect 27964 9546 27970 9610
rect 28034 9546 28186 9610
rect 27964 9540 28186 9546
rect 27966 8510 28186 9540
rect 28816 9488 34292 9708
rect 34512 9488 45822 9708
rect 28816 9444 45822 9488
rect 45522 8848 45822 9444
rect 27966 8504 28418 8510
rect 27966 8284 28192 8504
rect 28412 8284 28418 8504
rect 36281 8497 36527 8503
rect 28186 8278 28418 8284
rect 36255 8274 36281 8497
rect 36527 8274 37600 8491
rect 36568 8238 36791 8274
rect 19944 7372 20020 7378
rect 21449 7372 21696 7417
rect 19944 7308 19950 7372
rect 20014 7308 21696 7372
rect 19944 7302 20020 7308
rect 21623 7287 21696 7308
rect 33153 8015 36791 8238
rect 12533 6879 12753 6882
rect 10044 6815 12753 6879
rect 9980 6809 10044 6815
rect 10554 6716 10618 6722
rect 9894 6288 9958 6294
rect 10554 6288 10618 6652
rect 9958 6224 10618 6288
rect 9894 6218 9958 6224
rect 8748 5802 9818 5866
rect 12533 5864 12753 6815
rect 33153 6088 33376 8015
rect 37384 6938 37599 8274
rect 37384 6723 39365 6938
rect 33153 5877 33159 6088
rect 33370 5877 33376 6088
rect 33153 5865 33376 5877
rect 34286 6096 34518 6102
rect 5888 5620 5894 5672
rect 5946 5620 5952 5672
rect 7870 5694 7946 5700
rect 8748 5694 8812 5802
rect 9632 5799 9818 5802
rect 7870 5630 7876 5694
rect 7940 5630 8812 5694
rect 7870 5624 7946 5630
rect 5888 5608 5952 5620
rect 9757 5387 9818 5799
rect 11304 5858 11548 5864
rect 11304 5638 11316 5858
rect 11536 5638 11548 5858
rect 11304 5632 11548 5638
rect 12521 5858 12765 5864
rect 34286 5858 34518 5864
rect 12521 5638 12533 5858
rect 12756 5638 12765 5858
rect 12521 5632 12765 5638
rect 39150 5800 39365 6723
rect 48550 6422 48706 6486
rect 46959 6012 46965 6073
rect 47026 6012 47032 6073
rect 9750 5381 9824 5387
rect 9750 5320 9756 5381
rect 9818 5320 9824 5381
rect 9750 5314 9824 5320
rect 9711 4746 9786 4752
rect 9711 4687 9717 4746
rect 9780 4687 9786 4746
rect 9711 4681 9786 4687
rect 9719 4027 9778 4681
rect 9713 4021 9784 4027
rect 9713 3962 9719 4021
rect 9778 3962 9784 4021
rect 9713 3956 9784 3962
rect 9719 2741 9778 3956
rect 9713 2735 9784 2741
rect 9713 2676 9719 2735
rect 9778 2676 9784 2735
rect 9713 2670 9784 2676
rect 9719 1480 9778 2670
rect 11316 1488 11536 5632
rect 39150 5597 39156 5800
rect 39359 5597 39365 5800
rect 39150 5585 39365 5597
rect 9713 1474 9784 1480
rect 9713 1415 9719 1474
rect 9778 1415 9784 1474
rect 9713 1409 9784 1415
rect 11316 1280 11322 1488
rect 11530 1280 11536 1488
rect 11316 1268 11536 1280
rect 11939 1275 11998 1281
rect 13233 1277 13304 1288
rect 13233 1275 13239 1277
rect 11939 1269 13239 1275
rect 11939 1222 11945 1269
rect 11992 1222 13239 1269
rect 11939 1216 13239 1222
rect 11939 1210 11998 1216
rect 13233 1214 13239 1216
rect 13298 1276 13304 1277
rect 14518 1277 14590 1289
rect 15808 1277 15879 1283
rect 17094 1277 17165 1283
rect 18386 1277 18457 1283
rect 19674 1277 19745 1283
rect 20959 1277 21030 1283
rect 14518 1276 14524 1277
rect 13298 1217 14524 1276
rect 14584 1218 15814 1277
rect 15873 1218 17100 1277
rect 17159 1218 18392 1277
rect 18451 1218 19680 1277
rect 19739 1218 20965 1277
rect 21024 1218 21030 1277
rect 14584 1217 14590 1218
rect 13298 1214 13304 1217
rect 13233 1202 13304 1214
rect 14518 1205 14590 1217
rect 15808 1212 15879 1218
rect 17094 1212 17165 1218
rect 18386 1212 18457 1218
rect 19674 1212 19745 1218
rect 20959 1212 21030 1218
<< via1 >>
rect 27554 11426 27618 11490
rect 23821 11126 23894 11199
rect 9568 6815 9632 6879
rect 9370 6224 9434 6288
rect 7244 6036 7308 6100
rect 7700 6036 7764 6100
rect 10554 6988 10618 7056
rect 34292 9488 34512 9708
rect 36281 8274 36527 8497
rect 9980 6815 10044 6879
rect 10554 6652 10618 6716
rect 9894 6224 9958 6288
rect 34286 6090 34518 6096
rect 34286 5870 34292 6090
rect 34292 5870 34512 6090
rect 34512 5870 34518 6090
rect 34286 5864 34518 5870
rect 48960 6092 49036 6098
rect 46965 6067 47026 6073
rect 46965 6018 46971 6067
rect 46971 6018 47020 6067
rect 47020 6018 47026 6067
rect 46965 6012 47026 6018
rect 48960 6028 48966 6092
rect 48966 6028 49030 6092
rect 49030 6028 49036 6092
rect 48960 6022 49036 6028
rect 26382 -2357 26442 -2351
rect 26382 -2405 26388 -2357
rect 26388 -2405 26436 -2357
rect 26436 -2405 26442 -2357
rect 26382 -2411 26442 -2405
<< metal2 >>
rect 27554 11490 27618 11496
rect 27618 11426 29444 11490
rect 27554 11420 27618 11426
rect 23821 11199 23894 11205
rect 23821 11120 23894 11126
rect 29380 10074 29444 11426
rect 29380 10010 45994 10074
rect 34286 9488 34292 9708
rect 34512 9488 34518 9708
rect 10554 7056 10618 7062
rect 9562 6815 9568 6879
rect 9632 6815 9980 6879
rect 10044 6815 10050 6879
rect 10554 6716 10618 6988
rect 10548 6652 10554 6716
rect 10618 6652 10624 6716
rect 9370 6288 9434 6294
rect 9434 6224 9894 6288
rect 9958 6224 9964 6288
rect 9370 6218 9434 6224
rect 7700 6100 7764 6106
rect 7238 6036 7244 6100
rect 7308 6036 7700 6100
rect 34292 6096 34512 9488
rect 36293 9332 43589 9377
rect 45213 9332 45271 9336
rect 36293 9327 45276 9332
rect 36293 9269 45213 9327
rect 45271 9269 45276 9327
rect 36293 9264 45276 9269
rect 36293 9154 43589 9264
rect 45213 9260 45271 9264
rect 36293 8497 36516 9154
rect 45930 8634 45994 10010
rect 45500 8570 45994 8634
rect 46228 9332 46296 9341
rect 36275 8274 36281 8497
rect 36527 8274 36533 8497
rect 45500 6565 45564 8570
rect 46228 8434 46296 9264
rect 45656 8366 46296 8434
rect 45656 6664 45724 8366
rect 45656 6600 49030 6664
rect 45656 6598 45724 6600
rect 45500 6504 47026 6565
rect 45500 6502 45564 6504
rect 7700 6030 7764 6036
rect 46965 6073 47026 6504
rect 48966 6098 49030 6600
rect 46965 6006 47026 6012
<< via2 >>
rect 23821 11126 23894 11199
rect 45213 9269 45271 9327
rect 46228 9264 46296 9332
rect 26384 -2409 26440 -2353
<< metal3 >>
rect 46223 9332 46301 9337
rect 45208 9327 46228 9332
rect 45208 9269 45213 9327
rect 45271 9269 46228 9327
rect 45208 9264 46228 9269
rect 46296 9264 46301 9332
rect 46223 9259 46301 9264
rect 26379 -2349 26445 -2348
rect 26374 -2413 26380 -2349
rect 26444 -2413 26450 -2349
rect 26379 -2414 26445 -2413
<< via3 >>
rect 23816 11199 23899 11204
rect 23816 11126 23821 11199
rect 23821 11126 23894 11199
rect 23894 11126 23899 11199
rect 23816 11121 23899 11126
rect 26380 -2353 26444 -2349
rect 26380 -2409 26384 -2353
rect 26384 -2409 26440 -2353
rect 26440 -2409 26444 -2353
rect 26380 -2413 26444 -2409
<< metal4 >>
rect 26391 -2348 26432 -1945
rect 26379 -2349 26445 -2348
rect 26379 -2413 26380 -2349
rect 26444 -2413 26445 -2349
rect 26379 -2414 26445 -2413
<< via4 >>
rect 23698 11204 24018 11323
rect 23698 11121 23816 11204
rect 23816 11121 23899 11204
rect 23899 11121 24018 11204
rect 23698 11003 24018 11121
<< metal5 >>
rect 23674 11323 24042 11347
rect 23674 11003 23698 11323
rect 24018 11003 24042 11323
rect 23674 10979 24042 11003
use CNR_GR04_SSOPAMP  CNR_GR04_SSOPAMP_0
timestamp 1713446558
transform 1 0 5000 0 1 5200
box -5000 -5200 3412 3520
use CNR_GR04_SSOPAMP  CNR_GR04_SSOPAMP_1
timestamp 1713446558
transform 1 0 46090 0 1 5598
box -5000 -5200 3412 3520
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_1 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 26978 0 1 9412
box -184 -124 1528 1592
use CNRATR_PCH_8C4F0  CNRATR_PCH_8C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 11384 0 1 7224
box -184 -124 1912 1016
use CNRATR_PCH_8C4F0  CNRATR_PCH_8C4F0_1
timestamp 1695852000
transform 1 0 8984 0 1 7224
box -184 -124 1912 1016
use CNRATR_PCH_8C4F0  CNRATR_PCH_8C4F0_2
timestamp 1695852000
transform 1 0 19182 0 1 6898
box -184 -124 1912 1016
use sky130_fd_pr__cap_mim_m3_2_BESJ5K  sky130_fd_pr__cap_mim_m3_2_BESJ5K_0
timestamp 1713460579
transform 1 0 24159 0 1 4493
box -2349 -6600 2371 6600
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 3 1288 0 0 1288
timestamp 1705271942
transform 0 1 9100 -1 0 5704
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
array 0 7 1288 0 0 1288
timestamp 1705271942
transform 1 0 10993 0 1 500
box 0 0 1340 1340
use SUNTR_RPPO2  SUNTR_RPPO2_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1713272488
transform 1 0 37362 0 1 2154
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_1
timestamp 1713272488
transform 1 0 10700 0 1 2200
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_2
timestamp 1713272488
transform 1 0 32474 0 1 2432
box 0 0 2672 4236
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712309819
transform 0 -1 31850 1 0 400
box 0 0 8720 4236
<< labels >>
flabel locali 28036 10694 28100 10758 0 FreeSans 160 0 0 0 RESET
port 13 nsew
flabel locali 26805 8 45895 310 0 FreeSans 160 0 0 0 VSS
port 5 nsew
flabel metal1 48642 6422 48706 6486 0 FreeSans 160 0 0 0 COMPERATOR
port 27 nsew
flabel metal1 20904 11858 29116 12158 0 FreeSans 800 0 0 0 VDD_1V8
port 28 nsew
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713460579
<< metal4 >>
rect -2349 1039 2349 1080
rect -2349 561 2093 1039
rect 2329 561 2349 1039
rect -2349 520 2349 561
rect -2349 239 2349 280
rect -2349 -239 2093 239
rect 2329 -239 2349 239
rect -2349 -280 2349 -239
rect -2349 -561 2349 -520
rect -2349 -1039 2093 -561
rect 2329 -1039 2349 -561
rect -2349 -1080 2349 -1039
<< via4 >>
rect 2093 561 2329 1039
rect 2093 -239 2329 239
rect 2093 -1039 2329 -561
<< mimcap2 >>
rect -2269 960 1731 1000
rect -2269 640 -2229 960
rect 1691 640 1731 960
rect -2269 600 1731 640
rect -2269 160 1731 200
rect -2269 -160 -2229 160
rect 1691 -160 1731 160
rect -2269 -200 1731 -160
rect -2269 -640 1731 -600
rect -2269 -960 -2229 -640
rect 1691 -960 1731 -640
rect -2269 -1000 1731 -960
<< mimcap2contact >>
rect -2229 640 1691 960
rect -2229 -160 1691 160
rect -2229 -960 1691 -640
<< metal5 >>
rect -429 984 -109 1200
rect 2051 1039 2371 1200
rect -2253 960 1715 984
rect -2253 640 -2229 960
rect 1691 640 1715 960
rect -2253 616 1715 640
rect -429 184 -109 616
rect 2051 561 2093 1039
rect 2329 561 2371 1039
rect 2051 239 2371 561
rect -2253 160 1715 184
rect -2253 -160 -2229 160
rect 1691 -160 1715 160
rect -2253 -184 1715 -160
rect -429 -616 -109 -184
rect 2051 -239 2093 239
rect 2329 -239 2371 239
rect 2051 -561 2371 -239
rect -2253 -640 1715 -616
rect -2253 -960 -2229 -640
rect 1691 -960 1715 -640
rect -2253 -984 1715 -960
rect -429 -1200 -109 -984
rect 2051 -1039 2093 -561
rect 2329 -1039 2371 -561
rect 2051 -1200 2371 -1039
<< properties >>
string FIXED_BBOX -2349 520 1811 1080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20.00 l 2.00 val 88.36 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1712211083
<< error_p >>
rect -97 441 -33 447
rect 33 441 97 447
rect -97 407 -85 441
rect 33 407 45 441
rect -97 401 -33 407
rect 33 401 97 407
rect -97 -407 -33 -401
rect 33 -407 97 -401
rect -97 -441 -85 -407
rect 33 -441 45 -407
rect -97 -447 -33 -441
rect 33 -447 97 -441
<< nwell >>
rect -297 -579 297 579
<< pmos >>
rect -101 -360 -29 360
rect 29 -360 101 360
<< pdiff >>
rect -159 348 -101 360
rect -159 -348 -147 348
rect -113 -348 -101 348
rect -159 -360 -101 -348
rect -29 348 29 360
rect -29 -348 -17 348
rect 17 -348 29 348
rect -29 -360 29 -348
rect 101 348 159 360
rect 101 -348 113 348
rect 147 -348 159 348
rect 101 -360 159 -348
<< pdiffc >>
rect -147 -348 -113 348
rect -17 -348 17 348
rect 113 -348 147 348
<< nsubdiff >>
rect -261 509 -165 543
rect 165 509 261 543
rect -261 447 -227 509
rect 227 447 261 509
rect -261 -509 -227 -447
rect 227 -509 261 -447
rect -261 -543 -165 -509
rect 165 -543 261 -509
<< nsubdiffcont >>
rect -165 509 165 543
rect -261 -447 -227 447
rect 227 -447 261 447
rect -165 -543 165 -509
<< poly >>
rect -101 441 -29 457
rect -101 407 -85 441
rect -45 407 -29 441
rect -101 360 -29 407
rect 29 441 101 457
rect 29 407 45 441
rect 85 407 101 441
rect 29 360 101 407
rect -101 -407 -29 -360
rect -101 -441 -85 -407
rect -45 -441 -29 -407
rect -101 -457 -29 -441
rect 29 -407 101 -360
rect 29 -441 45 -407
rect 85 -441 101 -407
rect 29 -457 101 -441
<< polycont >>
rect -85 407 -45 441
rect 45 407 85 441
rect -85 -441 -45 -407
rect 45 -441 85 -407
<< locali >>
rect -261 509 -165 543
rect 165 509 261 543
rect -261 447 -227 509
rect 227 447 261 509
rect -101 407 -85 441
rect -45 407 -29 441
rect 29 407 45 441
rect 85 407 101 441
rect -147 348 -113 364
rect -147 -364 -113 -348
rect -17 348 17 364
rect -17 -364 17 -348
rect 113 348 147 364
rect 113 -364 147 -348
rect -101 -441 -85 -407
rect -45 -441 -29 -407
rect 29 -441 45 -407
rect 85 -441 101 -407
rect -261 -509 -227 -447
rect 227 -509 261 -447
rect -261 -543 -165 -509
rect 165 -543 261 -509
<< viali >>
rect -85 407 -45 441
rect 45 407 85 441
rect -147 -348 -113 348
rect -17 -348 17 348
rect 113 -348 147 348
rect -85 -441 -45 -407
rect 45 -441 85 -407
<< metal1 >>
rect -97 441 -33 447
rect -97 407 -85 441
rect -45 407 -33 441
rect -97 401 -33 407
rect 33 441 97 447
rect 33 407 45 441
rect 85 407 97 441
rect 33 401 97 407
rect -153 348 -107 360
rect -153 -348 -147 348
rect -113 -348 -107 348
rect -153 -360 -107 -348
rect -23 348 23 360
rect -23 -348 -17 348
rect 17 -348 23 348
rect -23 -360 23 -348
rect 107 348 153 360
rect 107 -348 113 348
rect 147 -348 153 348
rect 107 -360 153 -348
rect -97 -407 -33 -401
rect -97 -441 -85 -407
rect -45 -441 -33 -407
rect -97 -447 -33 -441
rect 33 -407 97 -401
rect 33 -441 45 -407
rect 85 -441 97 -407
rect 33 -447 97 -441
<< properties >>
string FIXED_BBOX -244 -526 244 526
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.6 l 0.36 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

.subckt top_verilog clk rst data_in start ready running d7 d6 d5 d4 d3 d2 d1 d0

adut [clk rst data_in start] [ready, running, d7 d6 d5 d4 d3 d2 d1 d0] null top 
.model top d_cosim simulation="./top.so" 
.ends
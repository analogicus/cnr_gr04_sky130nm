*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR04_DIFF-AMP_PK_lpe.spi
#else
.include ../../../work/xsch/CNR_GR04_DIFF-AMP_PK.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS     VSS     0       dc 0
VDD     VDD_1V8 0       dc 1.8
V_BIAS  IN_N    0       dc 0.9
V_IN    IN_P    IN_N    ac 1

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------



*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save ${VPORTS} all
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

set units = degrees
optran 0 0 0 1n 20u 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
*tran 10p 10n 1p
ac dec 20 1 1G
write
quit
#endif

.endc

.end

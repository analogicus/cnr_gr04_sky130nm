magic
tech sky130B
magscale 1 2
timestamp 1713440215
<< metal3 >>
rect -6798 2012 -2426 2040
rect -6798 -2012 -2510 2012
rect -2446 -2012 -2426 2012
rect -6798 -2040 -2426 -2012
rect -2186 2012 2186 2040
rect -2186 -2012 2102 2012
rect 2166 -2012 2186 2012
rect -2186 -2040 2186 -2012
rect 2426 2012 6798 2040
rect 2426 -2012 6714 2012
rect 6778 -2012 6798 2012
rect 2426 -2040 6798 -2012
<< via3 >>
rect -2510 -2012 -2446 2012
rect 2102 -2012 2166 2012
rect 6714 -2012 6778 2012
<< mimcap >>
rect -6758 1960 -2758 2000
rect -6758 -1960 -6718 1960
rect -2798 -1960 -2758 1960
rect -6758 -2000 -2758 -1960
rect -2146 1960 1854 2000
rect -2146 -1960 -2106 1960
rect 1814 -1960 1854 1960
rect -2146 -2000 1854 -1960
rect 2466 1960 6466 2000
rect 2466 -1960 2506 1960
rect 6426 -1960 6466 1960
rect 2466 -2000 6466 -1960
<< mimcapcontact >>
rect -6718 -1960 -2798 1960
rect -2106 -1960 1814 1960
rect 2506 -1960 6426 1960
<< metal4 >>
rect -2526 2012 -2430 2028
rect -6719 1960 -2797 1961
rect -6719 -1960 -6718 1960
rect -2798 -1960 -2797 1960
rect -6719 -1961 -2797 -1960
rect -2526 -2012 -2510 2012
rect -2446 -2012 -2430 2012
rect 2086 2012 2182 2028
rect -2107 1960 1815 1961
rect -2107 -1960 -2106 1960
rect 1814 -1960 1815 1960
rect -2107 -1961 1815 -1960
rect -2526 -2028 -2430 -2012
rect 2086 -2012 2102 2012
rect 2166 -2012 2182 2012
rect 6698 2012 6794 2028
rect 2505 1960 6427 1961
rect 2505 -1960 2506 1960
rect 6426 -1960 6427 1960
rect 2505 -1961 6427 -1960
rect 2086 -2028 2182 -2012
rect 6698 -2012 6714 2012
rect 6778 -2012 6794 2012
rect 6698 -2028 6794 -2012
<< properties >>
string FIXED_BBOX 2426 -2040 6506 2040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 20.00 l 20.00 val 815.2 carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713331242
<< error_p >>
rect -1202 160 -834 184
rect 296 160 664 184
rect -1202 -160 -1178 160
rect 296 -160 320 160
rect -1202 -184 -834 -160
rect 296 -184 664 -160
<< metal4 >>
rect -1298 239 -200 280
rect -1298 -239 -456 239
rect -220 -239 -200 239
rect -1298 -280 -200 -239
rect 200 239 1298 280
rect 200 -239 1042 239
rect 1278 -239 1298 239
rect 200 -280 1298 -239
<< via4 >>
rect -456 -239 -220 239
rect 1042 -239 1278 239
<< mimcap2 >>
rect -1218 160 -818 200
rect -1218 -160 -1178 160
rect -858 -160 -818 160
rect -1218 -200 -818 -160
rect 280 160 680 200
rect 280 -160 320 160
rect 640 -160 680 160
rect 280 -200 680 -160
<< mimcap2contact >>
rect -1178 -160 -858 160
rect 320 -160 640 160
<< metal5 >>
rect -498 239 -178 281
rect -1202 160 -834 184
rect -1202 -160 -1178 160
rect -858 -160 -834 160
rect -1202 -184 -834 -160
rect -498 -239 -456 239
rect -220 -239 -178 239
rect 1000 239 1320 281
rect 296 160 664 184
rect 296 -160 320 160
rect 640 -160 664 160
rect 296 -184 664 -160
rect -498 -281 -178 -239
rect 1000 -239 1042 239
rect 1278 -239 1320 239
rect 1000 -281 1320 -239
<< properties >>
string FIXED_BBOX 200 -280 760 280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

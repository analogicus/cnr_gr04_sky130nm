magic
tech sky130B
magscale 1 2
timestamp 1713446558
<< error_s >>
rect -4434 2684 -4428 2696
rect -4196 2684 -4190 2696
rect -4422 2672 -4410 2678
rect -4214 2672 -4202 2678
rect 1503 2642 1509 2654
rect 1607 2642 1613 2654
rect 1515 2630 1527 2636
rect 1589 2630 1601 2636
rect 876 2559 888 2565
rect 864 2541 870 2553
rect 864 2489 870 2501
rect 876 2477 888 2483
rect 1500 782 1518 788
rect 1580 782 1598 788
rect 1494 764 1500 782
rect 1598 764 1604 782
rect 1494 684 1500 702
rect 1598 684 1604 702
rect 1500 678 1518 684
rect 1580 678 1598 684
rect 448 498 454 510
rect 530 498 536 510
rect 460 486 472 492
rect 512 486 524 492
rect 1248 -1073 1254 -1061
rect 1330 -1073 1336 -1061
rect 1260 -1085 1272 -1079
rect 1312 -1085 1324 -1079
rect 1248 -2545 1254 -2533
rect 1330 -2545 1336 -2533
rect 1260 -2557 1272 -2551
rect 1312 -2557 1324 -2551
rect 704 -3314 716 -3308
rect 722 -3332 728 -3320
rect 722 -3384 728 -3372
rect 704 -3396 716 -3390
<< locali >>
rect -143 2642 1515 2728
rect 1601 2642 3243 2728
rect -155 690 1506 776
rect 1592 690 3255 776
rect -155 566 -69 690
rect 1185 585 1271 690
rect 1841 568 1927 690
rect 3169 547 3255 690
rect 876 430 1008 494
rect 2876 430 3012 494
rect -148 -800 1655 -714
rect -148 -934 -62 -800
rect 1569 -926 1655 -800
rect -165 -4449 -79 -4326
rect 1560 -4449 1646 -4335
rect -165 -4535 1646 -4449
rect 676 -4891 762 -4535
rect -497 -4952 3103 -4891
rect -497 -5026 1845 -4952
rect 1919 -5026 3103 -4952
rect -497 -5072 3103 -5026
rect -892 -5184 3103 -5072
rect -497 -5191 3103 -5184
<< viali >>
rect -4422 2684 -4202 2904
rect 1515 2642 1601 2728
rect 876 2489 940 2553
rect 2890 2495 2942 2547
rect 460 1922 524 1986
rect 882 1928 934 1980
rect 2460 1922 2524 1986
rect 1506 690 1592 776
rect 460 498 524 562
rect 2466 503 2518 555
rect 460 136 524 200
rect 2459 142 2511 194
rect 994 -1004 1046 -952
rect 1260 -1073 1324 -1009
rect -145 -1358 -93 -1306
rect 652 -1364 716 -1300
rect 1266 -1620 1318 -1568
rect 172 -1726 244 -1654
rect 927 -2452 979 -2400
rect 1260 -2545 1324 -2481
rect -119 -3378 -67 -3326
rect 652 -3384 716 -3320
rect -4320 -4455 -4260 -4395
rect 1845 -5026 1919 -4952
<< metal1 >>
rect -4422 3500 -345 3503
rect -4422 3283 3100 3500
rect -4422 2910 -4202 3283
rect -500 3200 3100 3283
rect -4428 2904 -4196 2910
rect -4428 2684 -4422 2904
rect -4202 2684 -4196 2904
rect 1515 2734 1601 3200
rect -4428 2678 -4196 2684
rect 1509 2728 1607 2734
rect 1509 2642 1515 2728
rect 1601 2642 1607 2728
rect 1509 2636 1607 2642
rect 870 2553 946 2559
rect 2884 2553 2948 2559
rect 870 2489 876 2553
rect 940 2547 2948 2553
rect 940 2495 2890 2547
rect 2942 2495 2948 2547
rect 940 2489 2948 2495
rect 870 2483 946 2489
rect 2884 2483 2948 2489
rect 454 1986 530 1998
rect 2448 1986 2536 1992
rect 454 1922 460 1986
rect 524 1980 946 1986
rect 524 1928 882 1980
rect 934 1928 946 1980
rect 524 1922 946 1928
rect 2448 1922 2460 1986
rect 2524 1922 2536 1986
rect 454 1910 530 1922
rect 2448 1916 2536 1922
rect 460 568 524 1910
rect 454 562 530 568
rect 454 498 460 562
rect 524 498 530 562
rect 454 492 530 498
rect 2460 555 2524 1916
rect 2460 503 2466 555
rect 2518 503 2524 555
rect 2460 491 2524 503
rect 454 200 530 212
rect 454 136 460 200
rect 524 194 2523 200
rect 524 142 2459 194
rect 2511 142 2523 194
rect 524 136 2523 142
rect 454 124 530 136
rect 1533 -530 1597 136
rect 1533 -594 1801 -530
rect 982 -952 1324 -946
rect 982 -1004 994 -952
rect 1046 -1003 1324 -952
rect 1046 -1004 1330 -1003
rect 982 -1009 1330 -1004
rect 982 -1010 1260 -1009
rect 1254 -1073 1260 -1010
rect 1324 -1073 1330 -1009
rect 1254 -1079 1330 -1073
rect -151 -1300 -87 -1294
rect 646 -1300 722 -1288
rect -151 -1306 652 -1300
rect -151 -1358 -145 -1306
rect -93 -1358 652 -1306
rect -151 -1364 652 -1358
rect 716 -1364 722 -1300
rect -151 -1370 -87 -1364
rect 646 -1376 722 -1364
rect 1260 -1568 1324 -1556
rect 1260 -1620 1266 -1568
rect 1318 -1620 1324 -1568
rect 160 -1654 256 -1648
rect 160 -1726 172 -1654
rect 244 -1726 256 -1654
rect 160 -1732 256 -1726
rect 172 -1877 244 -1732
rect -761 -1949 244 -1877
rect -4326 -4389 -4254 -4383
rect -761 -4389 -689 -1949
rect 915 -2191 921 -2127
rect 985 -2191 991 -2127
rect 921 -2400 985 -2191
rect 921 -2452 927 -2400
rect 979 -2452 985 -2400
rect 921 -2464 985 -2452
rect 1260 -2475 1324 -1620
rect 1737 -2127 1801 -594
rect 1534 -2191 1540 -2127
rect 1604 -2191 1801 -2127
rect 1254 -2481 1330 -2475
rect 1254 -2545 1260 -2481
rect 1324 -2545 1330 -2481
rect 1254 -2551 1330 -2545
rect 646 -3320 722 -3314
rect -131 -3326 652 -3320
rect -131 -3378 -119 -3326
rect -67 -3378 652 -3326
rect -131 -3384 652 -3378
rect 716 -3384 722 -3320
rect 646 -3390 722 -3384
rect -4326 -4395 -689 -4389
rect -4326 -4455 -4320 -4395
rect -4260 -4455 -689 -4395
rect -4326 -4461 -689 -4455
rect -4326 -4467 -4254 -4461
rect 1833 -5032 1839 -4946
rect 1925 -5032 1931 -4946
<< via1 >>
rect 1500 776 1598 782
rect 1500 690 1506 776
rect 1506 690 1592 776
rect 1592 690 1598 776
rect 1500 684 1598 690
rect 921 -2191 985 -2127
rect 1540 -2191 1604 -2127
rect 1839 -4952 1925 -4946
rect 1839 -5026 1845 -4952
rect 1845 -5026 1919 -4952
rect 1919 -5026 1925 -4952
rect 1839 -5032 1925 -5026
<< metal2 >>
rect 1506 494 1592 684
rect 1506 408 1713 494
rect 1627 -412 1713 408
rect 1627 -498 1925 -412
rect 921 -2127 985 -2121
rect 1540 -2127 1604 -2121
rect 985 -2191 1540 -2127
rect 921 -2197 985 -2191
rect 1540 -2197 1604 -2191
rect 1839 -4946 1925 -498
rect 1839 -5038 1925 -5032
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 1884 0 1 -276
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_1
timestamp 1695852000
transform 1 0 -116 0 1 -276
box -184 -124 1528 1016
use CNRATR_NCH_8C4F0  CNRATR_NCH_8C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -116 0 1 -1776
box -184 -124 1912 1016
use CNRATR_NCH_8C12F0  CNRATR_NCH_8C12F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -116 0 1 -4376
box -184 -124 1912 2168
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 1884 0 1 1224
box -184 -124 1528 1592
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_1
timestamp 1695852000
transform 1 0 -116 0 1 1224
box -184 -124 1528 1592
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712309819
transform 0 -1 -764 1 0 -5200
box 0 0 8720 4236
<< labels >>
flabel locali -497 -5191 1845 -4891 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 -500 3200 3100 3500 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel metal1 2460 555 2524 1922 0 FreeSans 1600 0 0 0 OPAMP_VOUT
port 5 nsew
flabel locali 942 430 1006 494 0 FreeSans 320 0 0 0 VIP
port 6 nsew
flabel locali 2948 430 3012 494 0 FreeSans 320 0 0 0 VIN
port 7 nsew
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713444105
<< error_s >>
rect -15375 -2260 -15369 -2248
rect -15271 -2260 -15265 -2248
rect -15363 -2272 -15351 -2266
rect -15289 -2272 -15277 -2266
rect -3743 -2296 -3737 -2216
rect -3663 -2296 -3657 -2216
rect -3743 -2302 -3657 -2296
rect -12024 -2408 -12012 -2402
rect -11520 -2412 -11514 -2406
rect -11462 -2412 -11456 -2406
rect -12036 -2426 -12030 -2414
rect -11526 -2416 -11520 -2412
rect -11456 -2416 -11450 -2412
rect 19085 -2460 19091 -2448
rect 19189 -2460 19195 -2448
rect -12036 -2478 -12030 -2466
rect 19097 -2472 19109 -2466
rect 19171 -2472 19183 -2466
rect -11526 -2476 -11520 -2472
rect -11456 -2476 -11450 -2472
rect -11520 -2482 -11514 -2476
rect -11462 -2482 -11456 -2476
rect -12024 -2490 -12012 -2484
rect 18476 -2602 18488 -2596
rect 18464 -2620 18470 -2608
rect 18464 -2672 18470 -2660
rect 18476 -2684 18488 -2678
rect -12440 -2696 -12428 -2690
rect -12388 -2696 -12376 -2690
rect -12452 -2714 -12446 -2702
rect -12370 -2714 -12364 -2702
rect -21106 -2770 -21100 -2758
rect -20868 -2770 -20862 -2758
rect -21094 -2782 -21082 -2776
rect -20886 -2782 -20874 -2776
rect -14440 -2908 -14428 -2902
rect -14388 -2908 -14376 -2902
rect -14452 -2926 -14446 -2914
rect -14370 -2926 -14364 -2914
rect 3066 -2930 3072 -2918
rect 3304 -2930 3310 -2918
rect 3078 -2942 3090 -2936
rect 3286 -2942 3298 -2936
rect 20060 -3108 20072 -3102
rect 20112 -3108 20124 -3102
rect 20048 -3126 20054 -3114
rect 20130 -3126 20136 -3114
rect -3759 -3237 -3753 -3235
rect -3695 -3237 -3689 -3235
rect -3759 -3241 -3745 -3237
rect -3703 -3241 -3689 -3237
rect -3765 -3246 -3683 -3241
rect -3765 -3247 -3754 -3246
rect -3763 -3250 -3754 -3247
rect -3750 -3247 -3744 -3246
rect -3704 -3247 -3698 -3246
rect -3750 -3250 -3698 -3247
rect -3694 -3247 -3683 -3246
rect -3694 -3250 -3685 -3247
rect -3763 -3255 -3685 -3250
rect -3759 -3256 -3692 -3255
rect -3759 -3296 -3754 -3256
rect -3750 -3259 -3698 -3256
rect -3750 -3293 -3741 -3259
rect -3750 -3296 -3698 -3293
rect -3759 -3297 -3692 -3296
rect -3763 -3302 -3685 -3297
rect -3763 -3305 -3754 -3302
rect -3765 -3306 -3754 -3305
rect -3750 -3305 -3698 -3302
rect -3750 -3306 -3744 -3305
rect -3704 -3306 -3698 -3305
rect -3694 -3305 -3685 -3302
rect -3694 -3306 -3683 -3305
rect -3765 -3311 -3683 -3306
rect -3759 -3315 -3745 -3311
rect -3703 -3315 -3689 -3311
rect -3759 -3317 -3753 -3315
rect -3695 -3317 -3689 -3315
rect -13905 -4321 -13893 -4315
rect -13831 -4321 -13819 -4315
rect -2807 -4327 -2801 -4321
rect -2739 -4327 -2733 -4321
rect -13917 -4339 -13911 -4327
rect -13813 -4339 -13807 -4327
rect -2813 -4332 -2727 -4327
rect -2813 -4333 -2802 -4332
rect -2733 -4333 -2727 -4332
rect -2807 -4395 -2802 -4333
rect -2813 -4396 -2802 -4395
rect -2733 -4396 -2727 -4395
rect -2813 -4401 -2727 -4396
rect -2807 -4407 -2801 -4401
rect -2739 -4407 -2733 -4401
rect -16452 -4606 -16446 -4594
rect -16370 -4606 -16364 -4594
rect -13263 -4612 -13257 -4606
rect -16440 -4618 -16428 -4612
rect -16388 -4618 -16376 -4612
rect -13256 -4618 -13251 -4612
rect -13256 -4673 -13251 -4668
rect -13324 -4674 -13318 -4673
rect -13257 -4674 -13251 -4673
rect -13318 -4680 -13312 -4674
rect -13263 -4680 -13257 -4674
rect -16440 -4894 -16428 -4888
rect -16452 -4912 -16446 -4900
rect -3456 -4952 -3450 -4940
rect -3374 -4952 -3368 -4940
rect -16452 -4964 -16446 -4952
rect -3444 -4964 -3432 -4958
rect -3392 -4964 -3380 -4958
rect -16440 -4976 -16428 -4970
rect -3866 -5448 -3860 -5442
rect -3796 -5448 -3790 -5442
rect -3872 -5454 -3866 -5448
rect -3790 -5454 -3784 -5448
rect -3872 -5524 -3866 -5518
rect -3790 -5524 -3784 -5518
rect -3866 -5530 -3860 -5524
rect -3796 -5530 -3790 -5524
rect -4397 -6252 -4340 -6243
rect -3188 -6252 -3143 -6243
rect -3757 -6271 -3739 -6265
rect -3677 -6271 -3659 -6265
rect -4397 -6286 -4306 -6277
rect -16248 -6292 -16236 -6286
rect -3763 -6289 -3757 -6271
rect -3659 -6289 -3653 -6271
rect -3222 -6286 -3143 -6277
rect -16260 -6310 -16254 -6298
rect -16260 -6362 -16254 -6350
rect -16248 -6374 -16236 -6368
rect -3763 -6369 -3757 -6351
rect -3659 -6369 -3653 -6351
rect -3757 -6375 -3739 -6369
rect -3677 -6375 -3659 -6369
rect -2476 -6454 -2475 -4310
rect 17523 -4623 17614 -4614
rect 18698 -4623 18797 -4614
rect 18883 -4623 18958 -4614
rect 19354 -4623 19437 -4614
rect 19523 -4623 19614 -4614
rect 20698 -4623 20777 -4614
rect 17523 -4657 17580 -4648
rect 18732 -4657 18797 -4648
rect 18883 -4657 18924 -4648
rect 19388 -4657 19437 -4648
rect 19523 -4657 19580 -4648
rect 20732 -4657 20777 -4648
rect 18048 -4806 18054 -4794
rect 18130 -4806 18136 -4794
rect 18470 -4808 18476 -4802
rect 18540 -4808 18546 -4802
rect 18060 -4818 18072 -4812
rect 18112 -4818 18124 -4812
rect 18464 -4814 18470 -4808
rect 18546 -4814 18552 -4808
rect 18464 -4884 18470 -4878
rect 18546 -4884 18552 -4878
rect 18470 -4890 18476 -4884
rect 18540 -4890 18546 -4884
rect 18060 -5088 18072 -5082
rect 20100 -5088 20112 -5082
rect 18048 -5106 18054 -5094
rect 20118 -5106 20124 -5094
rect 18048 -5158 18054 -5146
rect 20118 -5158 20124 -5146
rect 18060 -5170 18072 -5164
rect 20100 -5170 20112 -5164
rect 17523 -6023 17614 -6014
rect 19082 -6023 19157 -6014
rect 17523 -6057 17580 -6048
rect 19116 -6057 19157 -6048
rect 17516 -6482 17528 -6476
rect 17504 -6500 17510 -6488
rect -2701 -6601 -2695 -6595
rect -2633 -6601 -2627 -6595
rect -2707 -6606 -2621 -6601
rect -2707 -6607 -2696 -6606
rect -2627 -6607 -2621 -6606
rect -16734 -6648 -16716 -6642
rect -16668 -6648 -16650 -6642
rect -16740 -6666 -16734 -6648
rect -16650 -6666 -16644 -6648
rect -2701 -6669 -2696 -6607
rect -2707 -6670 -2696 -6669
rect -2627 -6670 -2621 -6669
rect -2707 -6675 -2621 -6670
rect -2701 -6681 -2695 -6675
rect -2633 -6681 -2627 -6675
rect -16740 -6732 -16734 -6714
rect -16650 -6732 -16644 -6714
rect -16734 -6738 -16716 -6732
rect -16668 -6738 -16650 -6732
rect -16977 -7363 -16906 -7362
rect -15438 -7363 -15343 -7362
rect -16977 -7397 -16940 -7396
rect -15404 -7397 -15343 -7396
rect -16082 -7482 -16076 -7476
rect -16012 -7482 -16006 -7476
rect -16088 -7488 -16082 -7482
rect -16006 -7488 -16000 -7482
rect -16088 -7558 -16082 -7552
rect -16006 -7558 -16000 -7552
rect -16082 -7564 -16076 -7558
rect -16012 -7564 -16006 -7558
rect -15660 -7562 -15659 -7556
rect -15597 -7562 -15596 -7556
rect -15672 -7580 -15666 -7568
rect -15590 -7580 -15584 -7568
rect -15672 -7632 -15666 -7620
rect -15590 -7632 -15584 -7620
rect -15660 -7644 -15648 -7638
rect -15608 -7644 -15596 -7638
rect -13740 -8616 -13730 -8582
rect -13702 -8649 -13692 -8588
rect -13014 -8647 -12991 -8588
rect -12976 -8616 -12953 -8582
rect -13637 -8649 -13631 -8647
rect -13655 -8661 -13643 -8655
rect -9580 -8816 -9570 -8782
rect -9542 -8830 -9532 -8768
rect -8288 -8816 -8282 -8782
rect -8250 -8828 -8244 -8769
rect -7566 -8827 -7551 -8768
rect -7528 -8816 -7513 -8782
rect -6278 -8820 -6257 -8773
rect -6240 -8816 -6219 -8782
rect -13744 -9621 -13620 -9615
rect -12496 -9621 -12372 -9615
rect -13710 -9655 -13654 -9649
rect -12462 -9655 -12406 -9649
rect -13014 -9749 -12991 -9732
rect -12976 -9787 -12953 -9770
rect -6313 -10040 -6301 -10034
rect -3344 -10038 -2795 -10037
rect -2476 -10038 -2475 -6502
rect 17504 -6552 17510 -6540
rect 17516 -6564 17528 -6558
rect 18860 -6782 18872 -6776
rect 18912 -6782 18924 -6776
rect 18848 -6800 18854 -6788
rect 18930 -6800 18936 -6788
rect 17778 -6848 17796 -6842
rect 17844 -6848 17862 -6842
rect 17772 -6866 17778 -6848
rect 17862 -6866 17868 -6848
rect 17772 -6932 17778 -6914
rect 17862 -6932 17868 -6914
rect 17778 -6938 17796 -6932
rect 17844 -6938 17862 -6932
rect 18438 -7682 18456 -7676
rect 18496 -7682 18514 -7676
rect 18432 -7700 18438 -7682
rect 18514 -7700 18520 -7682
rect 18432 -7758 18438 -7740
rect 18514 -7758 18520 -7740
rect 18438 -7764 18456 -7758
rect 18496 -7764 18514 -7758
rect -9588 -10104 -9570 -10070
rect -9550 -10106 -9532 -10045
rect -8308 -10104 -8282 -10070
rect -8270 -10107 -8244 -10046
rect -6325 -10047 -6319 -10046
rect -7008 -10104 -6994 -10070
rect -6970 -10108 -6956 -10047
rect -6325 -10110 -6319 -10108
rect -6278 -10110 -6252 -10046
rect -6240 -10104 -6214 -10070
rect -6313 -10122 -6301 -10116
rect -3344 -10357 -3343 -10038
rect -3024 -14867 -3023 -10357
rect -2637 -11528 -2158 -11492
rect -2637 -11812 -2539 -11528
rect -2514 -11549 -2508 -11547
rect -2286 -11549 -2280 -11547
rect -2514 -11552 -2500 -11549
rect -2294 -11552 -2280 -11549
rect -2514 -11553 -2491 -11552
rect -2520 -11558 -2514 -11553
rect -2509 -11558 -2491 -11553
rect -2303 -11553 -2280 -11552
rect -2303 -11558 -2285 -11553
rect -2280 -11558 -2274 -11553
rect -2520 -11559 -2509 -11558
rect -2518 -11567 -2509 -11559
rect -2515 -11576 -2509 -11567
rect -2285 -11559 -2274 -11558
rect -2285 -11567 -2276 -11559
rect -2285 -11576 -2279 -11567
rect -2515 -11773 -2509 -11764
rect -2518 -11781 -2509 -11773
rect -2520 -11782 -2509 -11781
rect -2285 -11773 -2279 -11764
rect -2285 -11781 -2276 -11773
rect -2285 -11782 -2274 -11781
rect -2520 -11787 -2514 -11782
rect -2509 -11787 -2491 -11782
rect -2514 -11788 -2491 -11787
rect -2303 -11787 -2285 -11782
rect -2280 -11787 -2274 -11782
rect -2303 -11788 -2280 -11787
rect -2514 -11791 -2500 -11788
rect -2294 -11791 -2280 -11788
rect -2514 -11793 -2508 -11791
rect -2286 -11793 -2280 -11791
rect -2255 -11812 -2158 -11528
rect -2317 -12400 -2158 -11812
rect -3024 -14868 -2483 -14867
rect -2798 -15187 -2483 -14868
rect -2262 -14880 -2163 -14548
rect -2478 -15200 -2163 -14880
rect -2262 -15507 -2163 -15200
<< locali >>
rect -15067 -2174 -13643 -2172
rect -17006 -2260 -15363 -2174
rect -15277 -2258 -13643 -2174
rect -15277 -2260 -15037 -2258
rect -13063 -2334 -11363 -2248
rect -11277 -2334 -9637 -2248
rect -4363 -2302 -3743 -2216
rect -3657 -2302 -3117 -2216
rect 17437 -2460 19097 -2374
rect 19183 -2460 20863 -2374
rect -17059 -4413 -13905 -4327
rect -13819 -4413 -13629 -4327
rect -17059 -4534 -16973 -4413
rect -15711 -4527 -15625 -4413
rect -15047 -4533 -14961 -4413
rect -13715 -4537 -13629 -4413
rect 17437 -4623 20753 -4537
rect 20839 -4623 20863 -4537
rect 17437 -4734 17523 -4623
rect 18797 -4723 18883 -4623
rect 19437 -4703 19523 -4623
rect 20777 -4743 20863 -4623
rect -17071 -5783 -15251 -5697
rect -17071 -5934 -16985 -5783
rect -15337 -5939 -15251 -5783
rect -16056 -6006 -15580 -5942
rect -15644 -6064 -15580 -6006
rect 17437 -6023 19243 -5937
rect 17437 -6134 17523 -6023
rect 19157 -6163 19243 -6023
rect -4483 -6277 -4397 -6166
rect -3143 -6277 -3057 -6177
rect -4483 -6363 -3751 -6277
rect -3665 -6363 -3057 -6277
rect -17063 -7363 -15257 -7277
rect -17063 -7483 -16977 -7363
rect -15343 -7482 -15257 -7363
rect 17437 -7543 19243 -7457
rect -10736 -7784 -10272 -7672
rect -7872 -7784 -7450 -7672
rect 17437 -7682 17523 -7543
rect 19157 -7703 19243 -7543
rect -13710 -9549 -13654 -9167
rect -12462 -9343 -12406 -9152
rect -12462 -9549 -12406 -9429
rect -13710 -9697 -13654 -9649
rect -12462 -9688 -12406 -9649
rect -13710 -9708 -13703 -9697
rect -13657 -9708 -13654 -9697
rect -17564 -11218 -17452 -10514
rect -13406 -11218 -13290 -10558
rect -10729 -11218 -10618 -7784
rect -10220 -8308 -10164 -8141
rect -8932 -8308 -8876 -8141
rect -7644 -8308 -7588 -8141
rect -6356 -8328 -6300 -8141
rect -10220 -9608 -10164 -9429
rect -8932 -9608 -8876 -9429
rect -7644 -9608 -7588 -9429
rect -6356 -9608 -6300 -9429
rect -2270 -10184 -1502 -9964
rect -7962 -11218 -7846 -10558
rect -3854 -10784 -2172 -10672
rect 6608 -10784 7146 -10672
rect 7578 -10782 7798 -9964
rect 11108 -10778 12386 -10666
rect -3854 -11218 -3742 -10784
rect 12274 -11218 12386 -10778
rect 12844 -11218 12956 -10716
rect -21792 -11249 12970 -11218
rect -21792 -11272 -14822 -11249
rect -21792 -11324 -15784 -11272
rect -15732 -11280 -14822 -11272
rect -15732 -11324 -15161 -11280
rect -21792 -11331 -15161 -11324
rect -15110 -11322 -14822 -11280
rect -14749 -11322 12970 -11249
rect -15110 -11331 12970 -11322
rect -21792 -11408 12970 -11331
rect -21792 -11460 -3854 -11408
rect -3802 -11451 12970 -11408
rect -3802 -11460 21291 -11451
rect -21792 -11499 21291 -11460
rect -21792 -11564 17231 -11499
rect -21792 -11776 -2503 -11564
rect -2291 -11573 17231 -11564
rect 17305 -11543 21291 -11499
rect 17305 -11573 19759 -11543
rect -2291 -11617 19759 -11573
rect 19833 -11617 21291 -11543
rect -2291 -11776 21291 -11617
rect -21792 -11810 21291 -11776
rect 11980 -12045 21291 -11810
rect 11980 -12284 12970 -12045
<< viali >>
rect -15363 -2260 -15277 -2174
rect -11363 -2334 -11277 -2248
rect -3743 -2302 -3657 -2216
rect -16024 -2432 -15960 -2368
rect -14020 -2426 -13968 -2374
rect -12024 -2478 -11960 -2414
rect -10024 -2420 -9960 -2414
rect -10024 -2472 -9954 -2420
rect -3518 -2472 -3466 -2420
rect 19097 -2460 19183 -2374
rect -10024 -2478 -9960 -2472
rect -21094 -2770 -20874 -2550
rect 18476 -2672 18540 -2608
rect 20474 -2666 20526 -2614
rect -12440 -2766 -12376 -2702
rect -10440 -2766 -10376 -2702
rect -1666 -2866 -1614 -2814
rect -16440 -2976 -16376 -2912
rect -16022 -2970 -15970 -2918
rect -14440 -2978 -14376 -2914
rect 3078 -2930 3298 -2710
rect 7605 -2915 7795 -2725
rect 13406 -2970 13626 -2750
rect 18066 -3116 18118 -3114
rect 18060 -3180 18124 -3116
rect 18494 -3174 18546 -3122
rect 20060 -3178 20124 -3114
rect -3741 -3293 -3707 -3259
rect -12534 -4314 -12466 -4246
rect -11432 -4262 -11380 -4210
rect -8560 -4242 -8508 -4190
rect -9714 -4314 -9646 -4246
rect -6934 -4294 -6866 -4226
rect -5690 -4248 -5638 -4196
rect -13905 -4413 -13819 -4327
rect -16440 -4606 -16376 -4542
rect -14434 -4604 -14382 -4552
rect -16022 -4666 -15970 -4614
rect -14018 -4667 -13969 -4618
rect 20753 -4623 20839 -4537
rect 18060 -4806 18124 -4742
rect 20066 -4802 20118 -4750
rect 18476 -4878 18540 -4814
rect 20476 -4878 20540 -4814
rect -16440 -4964 -16376 -4900
rect -14438 -4958 -14386 -4906
rect -3444 -4952 -3380 -4888
rect 18060 -5158 18124 -5094
rect 20048 -5158 20112 -5094
rect -3860 -5518 -3796 -5454
rect -3860 -6166 -3796 -6102
rect -16248 -6362 -16184 -6298
rect -15324 -6356 -15272 -6304
rect -3751 -6363 -3665 -6277
rect 17516 -6552 17580 -6488
rect 17914 -6546 17966 -6494
rect -15653 -6625 -15603 -6575
rect -16728 -6726 -16656 -6654
rect 18860 -6852 18924 -6788
rect 17784 -6926 17856 -6854
rect 17431 -7012 17517 -6926
rect -16076 -7552 -16012 -7488
rect -15660 -7632 -15596 -7568
rect 18444 -7752 18508 -7688
rect -16224 -8490 -16160 -8426
rect -15314 -8484 -15262 -8432
rect -13814 -8444 -13766 -8396
rect -13702 -8649 -13643 -8588
rect -13050 -8647 -12991 -8588
rect -20975 -9773 -20932 -9730
rect -13703 -9743 -13657 -9697
rect -13049 -9749 -12991 -9691
rect 18866 -7826 18918 -7774
rect 17514 -8684 17566 -8632
rect 18252 -8690 18316 -8626
rect -9542 -8830 -9483 -8768
rect -8250 -8828 -8191 -8769
rect -7610 -8827 -7551 -8768
rect -6304 -8820 -6257 -8773
rect 17423 -9712 17509 -9626
rect -9550 -10106 -9489 -10045
rect -8270 -10107 -8209 -10046
rect -6970 -10108 -6909 -10047
rect -6313 -10110 -6252 -10046
rect 3078 -10184 3298 -9964
rect 13510 -10130 13570 -10070
rect -15784 -11324 -15732 -11272
rect -15161 -11331 -15110 -11280
rect -14822 -11322 -14749 -11249
rect -3854 -11460 -3802 -11408
rect -2503 -11776 -2291 -11564
rect 17231 -11573 17305 -11499
rect 19759 -11617 19833 -11543
<< metal1 >>
rect -19760 -1250 19410 -1240
rect -21094 -1470 19410 -1250
rect -21094 -2544 -20874 -1470
rect -19760 -1540 19410 -1470
rect -15363 -2168 -15277 -1540
rect -15369 -2174 -15271 -2168
rect -15369 -2260 -15363 -2174
rect -15277 -2260 -15271 -2174
rect -11363 -2236 -11277 -1540
rect -3743 -2216 -3657 -1540
rect -15369 -2266 -15271 -2260
rect -11369 -2248 -11271 -2236
rect -11369 -2334 -11363 -2248
rect -11277 -2334 -11271 -2248
rect -11369 -2346 -11271 -2334
rect -16030 -2368 -15954 -2356
rect -14026 -2368 -13962 -2362
rect -16030 -2432 -16024 -2368
rect -15960 -2374 -13962 -2368
rect -15960 -2426 -14020 -2374
rect -13968 -2426 -13962 -2374
rect -15960 -2432 -13962 -2426
rect -16030 -2444 -15954 -2432
rect -14026 -2438 -13962 -2432
rect -12030 -2414 -11954 -2408
rect -12030 -2478 -12024 -2414
rect -11960 -2476 -11520 -2414
rect -10036 -2414 -9948 -2408
rect -11456 -2476 -10024 -2414
rect -9960 -2420 -3454 -2414
rect -9954 -2472 -3518 -2420
rect -3466 -2472 -3454 -2420
rect -11960 -2478 -10024 -2476
rect -9960 -2478 -3454 -2472
rect -12030 -2484 -11954 -2478
rect -10036 -2484 -9948 -2478
rect -21100 -2550 -20868 -2544
rect -21100 -2770 -21094 -2550
rect -20874 -2770 -20868 -2550
rect -21100 -2776 -20868 -2770
rect -12446 -2702 -12370 -2696
rect -12446 -2766 -12440 -2702
rect -12376 -2766 -12370 -2702
rect -12446 -2772 -12370 -2766
rect -10452 -2702 -10364 -2696
rect -10452 -2766 -10440 -2702
rect -10376 -2766 -10364 -2702
rect 3078 -2704 3298 -1540
rect 13406 -1846 13626 -1540
rect 6840 -1910 17274 -1846
rect -10452 -2772 -10364 -2766
rect 3072 -2710 3304 -2704
rect -16446 -2912 -16370 -2900
rect -16446 -2976 -16440 -2912
rect -16376 -2918 -15958 -2912
rect -16376 -2970 -16022 -2918
rect -15970 -2970 -15958 -2918
rect -16376 -2976 -15958 -2970
rect -14446 -2914 -14370 -2908
rect -16446 -2988 -16370 -2976
rect -14446 -2978 -14440 -2914
rect -14376 -2978 -14370 -2914
rect -14446 -2984 -14370 -2978
rect -16440 -4536 -16376 -2988
rect -14440 -3788 -14376 -2984
rect -12440 -3284 -12376 -2772
rect -13320 -3348 -12376 -3284
rect -13472 -3480 -13466 -3416
rect -13402 -3480 -13396 -3416
rect -14644 -4024 -14580 -4018
rect -16028 -4088 -14644 -4024
rect -16446 -4542 -16370 -4536
rect -16446 -4606 -16440 -4542
rect -16376 -4606 -16370 -4542
rect -16446 -4612 -16370 -4606
rect -16028 -4614 -15964 -4088
rect -14644 -4094 -14580 -4088
rect -16028 -4666 -16022 -4614
rect -15970 -4666 -15964 -4614
rect -14440 -4552 -14376 -3852
rect -13466 -4024 -13402 -3480
rect -14188 -4088 -14182 -4024
rect -14118 -4088 -13402 -4024
rect -13911 -4327 -13813 -4321
rect -13911 -4413 -13905 -4327
rect -13819 -4413 -13813 -4327
rect -13911 -4419 -13813 -4413
rect -14440 -4604 -14434 -4552
rect -14382 -4604 -14376 -4552
rect -14440 -4616 -14376 -4604
rect -14024 -4612 -13963 -4606
rect -16028 -4678 -15964 -4666
rect -14024 -4679 -13963 -4673
rect -16446 -4900 -16370 -4894
rect -16446 -4964 -16440 -4900
rect -16376 -4906 -14374 -4900
rect -16376 -4908 -14438 -4906
rect -16376 -4964 -15352 -4908
rect -16446 -4970 -16370 -4964
rect -15358 -4973 -15352 -4964
rect -15287 -4958 -14438 -4908
rect -14386 -4958 -14374 -4906
rect -15287 -4964 -14374 -4958
rect -15287 -4973 -15281 -4964
rect -13905 -5481 -13819 -4419
rect -14829 -5567 -13819 -5481
rect -13318 -4612 -13257 -3348
rect -13124 -3416 -13060 -3410
rect -10440 -3414 -10376 -2772
rect -2512 -2808 -2448 -2806
rect -1672 -2808 -1608 -2802
rect -2512 -2814 -1608 -2808
rect -2512 -2866 -1666 -2814
rect -1614 -2866 -1608 -2814
rect -2512 -2872 -1608 -2866
rect -3747 -3250 -3701 -3247
rect -3747 -3305 -3701 -3302
rect -10440 -3416 -5632 -3414
rect -13060 -3478 -5632 -3416
rect -13060 -3480 -10376 -3478
rect -13124 -3486 -13060 -3480
rect -11438 -4210 -11374 -3480
rect -16254 -6298 -16178 -6292
rect -16254 -6362 -16248 -6298
rect -16184 -6304 -15260 -6298
rect -16184 -6356 -15324 -6304
rect -15272 -6356 -15260 -6304
rect -16184 -6362 -15260 -6356
rect -16254 -6368 -16178 -6362
rect -15665 -6575 -15591 -6569
rect -15665 -6625 -15653 -6575
rect -15603 -6625 -15591 -6575
rect -15665 -6631 -15591 -6625
rect -16088 -7558 -16082 -7482
rect -16006 -7558 -16000 -7482
rect -15659 -7562 -15597 -6631
rect -15492 -7184 -15428 -6362
rect -15492 -7248 -15104 -7184
rect -15666 -7568 -15590 -7562
rect -15666 -7632 -15660 -7568
rect -15596 -7632 -15590 -7568
rect -15666 -7638 -15590 -7632
rect -16230 -8426 -16154 -8414
rect -16230 -8490 -16224 -8426
rect -16160 -8432 -15250 -8426
rect -16160 -8484 -15314 -8432
rect -15262 -8484 -15250 -8432
rect -16160 -8490 -15250 -8484
rect -16230 -8502 -16154 -8490
rect -20981 -9724 -20926 -9718
rect -20981 -9785 -20926 -9779
rect -15790 -11272 -15726 -8490
rect -15790 -11324 -15784 -11272
rect -15732 -11324 -15726 -11272
rect -15790 -11336 -15726 -11324
rect -15167 -11280 -15104 -7248
rect -15167 -11331 -15161 -11280
rect -15110 -11331 -15104 -11280
rect -15167 -11343 -15104 -11331
rect -14828 -11249 -14743 -5567
rect -13318 -7865 -13257 -4674
rect -13820 -7925 -13257 -7865
rect -13820 -8396 -13760 -7925
rect -13318 -7926 -13257 -7925
rect -12540 -4246 -12460 -4234
rect -12540 -4314 -12534 -4246
rect -12466 -4314 -12460 -4246
rect -11438 -4262 -11432 -4210
rect -11380 -4262 -11374 -4210
rect -8566 -4190 -8502 -3478
rect -11438 -4274 -11374 -4262
rect -9726 -4246 -9634 -4240
rect -12540 -7920 -12460 -4314
rect -9726 -4314 -9714 -4246
rect -9646 -4314 -9634 -4246
rect -8566 -4242 -8560 -4190
rect -8508 -4242 -8502 -4190
rect -5696 -4196 -5632 -3478
rect -8566 -4254 -8502 -4242
rect -6940 -4226 -6860 -4214
rect -9726 -4320 -9634 -4314
rect -6940 -4294 -6934 -4226
rect -6866 -4294 -6860 -4226
rect -5696 -4248 -5690 -4196
rect -5638 -4248 -5632 -4196
rect -5696 -4260 -5632 -4248
rect -9720 -7920 -9640 -4320
rect -6940 -7920 -6860 -4294
rect -2512 -4468 -2448 -2872
rect -1672 -2878 -1608 -2872
rect 3072 -2930 3078 -2710
rect 3298 -2930 3304 -2710
rect 6840 -2719 6904 -1910
rect 3072 -2936 3304 -2930
rect 6739 -2725 7807 -2719
rect 6739 -2915 7605 -2725
rect 7795 -2915 7807 -2725
rect 13406 -2738 13626 -1910
rect 6739 -2921 7807 -2915
rect 13400 -2750 13632 -2738
rect -3444 -4530 -2448 -4468
rect -3444 -4532 -2512 -4530
rect -3444 -4882 -3380 -4532
rect -3450 -4888 -3374 -4882
rect -3450 -4952 -3444 -4888
rect -3380 -4952 -3374 -4888
rect -3450 -4958 -3374 -4952
rect -3872 -5524 -3866 -5448
rect -3790 -5524 -3784 -5448
rect -3872 -6102 -3784 -6096
rect -3872 -6166 -3860 -6102
rect -3796 -6166 -3784 -6102
rect -3872 -6172 -3784 -6166
rect -3860 -6606 -3796 -6172
rect -3860 -6670 -2696 -6606
rect -2632 -6670 -2626 -6606
rect -12540 -8000 -5340 -7920
rect -13820 -8444 -13814 -8396
rect -13766 -8444 -13760 -8396
rect -13820 -8456 -13760 -8444
rect -13708 -8588 -13637 -8582
rect -13062 -8588 -12979 -8582
rect -13708 -8649 -13702 -8588
rect -13643 -8647 -13050 -8588
rect -12991 -8647 -12979 -8588
rect -13643 -8649 -13637 -8647
rect -13708 -8655 -13637 -8649
rect -13062 -8653 -12979 -8647
rect -13049 -9685 -12991 -8653
rect -9541 -8756 -9482 -8000
rect -9548 -8762 -9477 -8756
rect -9554 -8768 -9471 -8762
rect -9554 -8830 -9542 -8768
rect -9483 -8769 -9471 -8768
rect -8256 -8768 -8185 -8757
rect -7616 -8767 -7545 -8762
rect -7616 -8768 -6245 -8767
rect -8256 -8769 -7610 -8768
rect -9483 -8828 -8250 -8769
rect -8191 -8827 -7610 -8769
rect -7551 -8773 -6245 -8768
rect -7551 -8820 -6304 -8773
rect -6257 -8820 -6245 -8773
rect -7551 -8826 -6245 -8820
rect -7551 -8827 -7545 -8826
rect -8191 -8828 -8185 -8827
rect -9483 -8830 -9471 -8828
rect -9554 -8833 -9471 -8830
rect -9549 -8842 -9477 -8833
rect -8256 -8840 -8185 -8828
rect -7616 -8833 -7545 -8827
rect -13055 -9691 -12985 -9685
rect -13715 -9697 -13049 -9691
rect -13715 -9743 -13703 -9697
rect -13657 -9743 -13049 -9697
rect -13715 -9749 -13049 -9743
rect -12991 -9749 -12985 -9691
rect -13055 -9755 -12985 -9749
rect -9549 -10039 -9488 -8842
rect 3072 -9964 3304 -9952
rect 6739 -9964 6941 -2921
rect 13400 -2970 13406 -2750
rect 13626 -2970 13632 -2750
rect 13400 -2982 13632 -2970
rect 17210 -4106 17274 -1910
rect 19097 -2368 19183 -1540
rect 19091 -2374 19189 -2368
rect 19091 -2460 19097 -2374
rect 19183 -2460 19189 -2374
rect 19091 -2466 19189 -2460
rect 18470 -2608 18546 -2602
rect 18470 -2672 18476 -2608
rect 18540 -2614 20538 -2608
rect 18540 -2666 20474 -2614
rect 20526 -2666 20538 -2614
rect 18540 -2672 20538 -2666
rect 18470 -2678 18546 -2672
rect 18060 -3110 18124 -3102
rect 18054 -3114 18130 -3110
rect 18054 -3116 18066 -3114
rect 18118 -3116 18130 -3114
rect 20054 -3114 20130 -3108
rect 18054 -3180 18060 -3116
rect 18124 -3122 18558 -3116
rect 18124 -3174 18494 -3122
rect 18546 -3174 18558 -3122
rect 18124 -3180 18558 -3174
rect 20054 -3178 20060 -3114
rect 20124 -3178 20130 -3114
rect 18054 -3186 18130 -3180
rect 20054 -3184 20130 -3178
rect 17578 -4106 17642 -4100
rect 17210 -4170 17578 -4106
rect 17578 -4176 17642 -4170
rect 18060 -4736 18124 -3186
rect 18054 -4742 18130 -4736
rect 18054 -4806 18060 -4742
rect 18124 -4806 18130 -4742
rect 18054 -4812 18130 -4806
rect 20060 -4750 20124 -3184
rect 20747 -4537 20845 -4525
rect 20747 -4623 20753 -4537
rect 20839 -4623 21133 -4537
rect 20747 -4635 20845 -4623
rect 20060 -4802 20066 -4750
rect 20118 -4802 20124 -4750
rect 18464 -4884 18470 -4808
rect 18546 -4884 18552 -4808
rect 20060 -4814 20124 -4802
rect 20464 -4814 20552 -4808
rect 20464 -4820 20476 -4814
rect 20540 -4820 20552 -4814
rect 20464 -4884 20470 -4820
rect 20546 -4884 20552 -4820
rect 20470 -4890 20546 -4884
rect 18054 -5094 18130 -5088
rect 19102 -5094 19108 -5088
rect 18054 -5158 18060 -5094
rect 18124 -5152 19108 -5094
rect 19172 -5094 19178 -5088
rect 20042 -5094 20118 -5088
rect 19172 -5152 20048 -5094
rect 18124 -5158 20048 -5152
rect 20112 -5158 20118 -5094
rect 18054 -5164 18130 -5158
rect 20042 -5164 20118 -5158
rect 21047 -5865 21133 -4623
rect 19753 -5951 21133 -5865
rect 17510 -6488 17586 -6482
rect 17510 -6552 17516 -6488
rect 17580 -6494 17978 -6488
rect 17580 -6546 17914 -6494
rect 17966 -6546 17978 -6494
rect 17580 -6552 17978 -6546
rect 17510 -6558 17586 -6552
rect 18854 -6788 18930 -6782
rect 17419 -6926 17529 -6920
rect 17419 -7012 17431 -6926
rect 17517 -7012 17529 -6926
rect 18854 -6852 18860 -6788
rect 18924 -6852 18930 -6788
rect 18854 -6858 18930 -6852
rect 17419 -7018 17529 -7012
rect 17431 -7175 17517 -7018
rect 17225 -7261 17517 -7175
rect 17225 -9825 17311 -7261
rect 18860 -7774 18924 -6858
rect 18860 -7826 18866 -7774
rect 18918 -7826 18924 -7774
rect 18860 -7838 18924 -7826
rect 18246 -8626 18322 -8614
rect 17502 -8632 18252 -8626
rect 17502 -8684 17514 -8632
rect 17566 -8684 18252 -8632
rect 17502 -8690 18252 -8684
rect 18316 -8690 18322 -8626
rect 18246 -8702 18322 -8690
rect 17411 -9626 17521 -9620
rect 17411 -9712 17423 -9626
rect 17509 -9712 17521 -9626
rect 17411 -9718 17521 -9712
rect 17423 -9825 17509 -9718
rect 17225 -9911 17509 -9825
rect -9556 -10045 -9483 -10039
rect -8276 -10045 -8203 -10040
rect -9556 -10106 -9550 -10045
rect -9489 -10046 -8203 -10045
rect -6976 -10046 -6903 -10035
rect -9489 -10106 -8270 -10046
rect -9556 -10112 -9483 -10106
rect -8276 -10107 -8270 -10106
rect -8209 -10047 -6903 -10046
rect -6319 -10046 -6246 -10040
rect -6319 -10047 -6313 -10046
rect -8209 -10107 -6970 -10047
rect -8276 -10113 -8203 -10107
rect -6976 -10108 -6970 -10107
rect -6909 -10108 -6313 -10047
rect -6976 -10120 -6903 -10108
rect -6319 -10110 -6313 -10108
rect -6252 -10110 -6246 -10046
rect -6319 -10116 -6246 -10110
rect 3072 -10184 3078 -9964
rect 3298 -10184 6950 -9964
rect 13504 -10064 13576 -10058
rect 13504 -10142 13576 -10136
rect 3072 -10196 3304 -10184
rect -14828 -11322 -14822 -11249
rect -14749 -11322 -14743 -11249
rect -14828 -11334 -14743 -11322
rect -3866 -11466 -3860 -11402
rect -3796 -11466 -3790 -11402
rect 17225 -11499 17311 -9911
rect 17225 -11573 17231 -11499
rect 17305 -11573 17311 -11499
rect 19753 -11537 19839 -5951
rect 17225 -11585 17311 -11573
rect 19747 -11543 19845 -11537
rect 19747 -11617 19759 -11543
rect 19833 -11617 19845 -11543
rect 19747 -11623 19845 -11617
<< via1 >>
rect -11520 -2476 -11456 -2412
rect -13466 -3480 -13402 -3416
rect -14440 -3852 -14376 -3788
rect -14644 -4088 -14580 -4024
rect -14182 -4088 -14118 -4024
rect -14024 -4618 -13963 -4612
rect -14024 -4667 -14018 -4618
rect -14018 -4667 -13969 -4618
rect -13969 -4667 -13963 -4618
rect -14024 -4673 -13963 -4667
rect -15352 -4973 -15287 -4908
rect -3750 -3259 -3698 -3250
rect -3750 -3293 -3741 -3259
rect -3741 -3293 -3707 -3259
rect -3707 -3293 -3698 -3259
rect -3750 -3302 -3698 -3293
rect -13124 -3480 -13060 -3416
rect -13318 -4674 -13257 -4612
rect -16734 -6654 -16650 -6648
rect -16734 -6726 -16728 -6654
rect -16728 -6726 -16656 -6654
rect -16656 -6726 -16650 -6654
rect -16734 -6732 -16650 -6726
rect -16082 -7488 -16006 -7482
rect -16082 -7552 -16076 -7488
rect -16076 -7552 -16012 -7488
rect -16012 -7552 -16006 -7488
rect -16082 -7558 -16006 -7552
rect -20981 -9730 -20926 -9724
rect -20981 -9773 -20975 -9730
rect -20975 -9773 -20932 -9730
rect -20932 -9773 -20926 -9730
rect -20981 -9779 -20926 -9773
rect -3866 -5454 -3790 -5448
rect -3866 -5518 -3860 -5454
rect -3860 -5518 -3796 -5454
rect -3796 -5518 -3790 -5454
rect -3866 -5524 -3790 -5518
rect -3757 -6277 -3659 -6271
rect -3757 -6363 -3751 -6277
rect -3751 -6363 -3665 -6277
rect -3665 -6363 -3659 -6277
rect -3757 -6369 -3659 -6363
rect -2696 -6670 -2632 -6606
rect 17578 -4170 17642 -4106
rect 18470 -4814 18546 -4808
rect 18470 -4878 18476 -4814
rect 18476 -4878 18540 -4814
rect 18540 -4878 18546 -4814
rect 18470 -4884 18546 -4878
rect 20470 -4878 20476 -4820
rect 20476 -4878 20540 -4820
rect 20540 -4878 20546 -4820
rect 20470 -4884 20546 -4878
rect 19108 -5152 19172 -5088
rect 17778 -6854 17862 -6848
rect 17778 -6926 17784 -6854
rect 17784 -6926 17856 -6854
rect 17856 -6926 17862 -6854
rect 17778 -6932 17862 -6926
rect 18438 -7688 18514 -7682
rect 18438 -7752 18444 -7688
rect 18444 -7752 18508 -7688
rect 18508 -7752 18514 -7688
rect 18438 -7758 18514 -7752
rect 13504 -10070 13576 -10064
rect 13504 -10130 13510 -10070
rect 13510 -10130 13570 -10070
rect 13570 -10130 13576 -10070
rect 13504 -10136 13576 -10130
rect -3860 -11408 -3796 -11402
rect -3860 -11460 -3854 -11408
rect -3854 -11460 -3802 -11408
rect -3802 -11460 -3796 -11408
rect -3860 -11466 -3796 -11460
rect -2509 -11564 -2285 -11558
rect -2509 -11776 -2503 -11564
rect -2503 -11776 -2291 -11564
rect -2291 -11776 -2285 -11564
rect -2509 -11782 -2285 -11776
<< metal2 >>
rect -2802 -2006 17208 -1942
rect -11525 -2472 -11520 -2416
rect -11456 -2472 -11451 -2416
rect -13466 -3416 -13402 -3410
rect -13402 -3480 -13124 -3416
rect -13060 -3480 -13054 -3416
rect -13466 -3486 -13402 -3480
rect -14449 -3852 -14440 -3788
rect -14376 -3852 -14367 -3788
rect -14182 -4024 -14118 -4018
rect -14650 -4088 -14644 -4024
rect -14580 -4088 -14182 -4024
rect -14182 -4094 -14118 -4088
rect -2802 -4332 -2738 -2006
rect 17144 -4248 17208 -2006
rect 17572 -4170 17578 -4106
rect 17642 -4170 20540 -4106
rect 17144 -4312 18540 -4248
rect -2802 -4405 -2738 -4396
rect -14030 -4673 -14024 -4612
rect -13963 -4673 -13318 -4612
rect -13257 -4673 -13256 -4612
rect 18476 -4808 18540 -4312
rect 20476 -4820 20540 -4170
rect 20464 -4884 20470 -4820
rect 20546 -4884 20552 -4820
rect -15352 -4908 -15287 -4902
rect -15352 -5528 -15287 -4973
rect 19108 -5088 19172 -5082
rect -15352 -5593 -15007 -5528
rect -16728 -6898 -16656 -6732
rect -17396 -6970 -16656 -6898
rect -17387 -9724 -17332 -6970
rect -15072 -7028 -15007 -5593
rect -3860 -6277 -3796 -5524
rect 19108 -5748 19172 -5152
rect 19108 -5812 19532 -5748
rect -3865 -6363 -3757 -6277
rect -16076 -7092 -15007 -7028
rect -16076 -7482 -16012 -7092
rect -20987 -9779 -20981 -9724
rect -20926 -9779 -17332 -9724
rect -3860 -11402 -3796 -6363
rect -2696 -6606 -2632 -6597
rect -2696 -6679 -2632 -6670
rect 17784 -7044 17856 -6932
rect 17124 -7116 17856 -7044
rect 17124 -10064 17196 -7116
rect 19468 -7188 19532 -5812
rect 18444 -7252 19532 -7188
rect 18444 -7682 18508 -7252
rect 13498 -10136 13504 -10064
rect 13576 -10136 17196 -10064
rect -3860 -11472 -3796 -11466
<< via2 >>
rect -11516 -2472 -11460 -2416
rect -3754 -3250 -3694 -3246
rect -3754 -3302 -3750 -3250
rect -3750 -3302 -3698 -3250
rect -3698 -3302 -3694 -3250
rect -3754 -3306 -3694 -3302
rect -14440 -3852 -14376 -3788
rect -2802 -4396 -2738 -4332
rect -2696 -6670 -2632 -6606
rect -2509 -11782 -2285 -11558
<< metal3 >>
rect -11521 -2416 -11455 -2411
rect -11521 -2472 -11516 -2416
rect -11460 -2472 -11455 -2416
rect -11521 -2477 -11455 -2472
rect -11520 -3514 -11456 -2477
rect -13242 -3578 -11456 -3514
rect -14445 -3788 -14371 -3783
rect -13242 -3788 -13178 -3578
rect -14445 -3852 -14440 -3788
rect -14376 -3852 -13178 -3788
rect -14445 -3857 -14371 -3852
<< via3 >>
rect -3759 -3246 -3689 -3241
rect -3759 -3306 -3754 -3246
rect -3754 -3306 -3694 -3246
rect -3694 -3306 -3689 -3246
rect -3759 -3311 -3689 -3306
rect -2807 -4332 -2733 -4327
rect -2807 -4396 -2802 -4332
rect -2802 -4396 -2738 -4332
rect -2738 -4396 -2733 -4332
rect -2807 -4401 -2733 -4396
rect -2701 -6606 -2627 -6601
rect -2701 -6670 -2696 -6606
rect -2696 -6670 -2632 -6606
rect -2632 -6670 -2627 -6606
rect -2701 -6675 -2627 -6670
rect -2514 -11558 -2280 -11553
rect -2514 -11782 -2509 -11558
rect -2509 -11782 -2285 -11558
rect -2285 -11782 -2280 -11558
rect -2514 -11787 -2280 -11782
<< via4 >>
rect -3884 -3241 -3564 -3116
rect -3884 -3311 -3759 -3241
rect -3759 -3311 -3689 -3241
rect -3689 -3311 -3564 -3241
rect -3884 -3436 -3564 -3311
rect -2930 -4327 -2610 -4204
rect -2930 -4334 -2807 -4327
rect -2946 -4401 -2807 -4334
rect -2807 -4401 -2733 -4327
rect -2733 -4401 -2610 -4327
rect -2946 -4524 -2610 -4401
rect -2946 -4606 -2674 -4524
rect -2824 -6601 -2504 -6478
rect -2824 -6675 -2701 -6601
rect -2701 -6675 -2627 -6601
rect -2627 -6675 -2504 -6601
rect -2824 -6798 -2504 -6675
rect -2515 -11553 -2279 -11552
rect -2515 -11787 -2514 -11553
rect -2514 -11787 -2280 -11553
rect -2280 -11787 -2279 -11553
rect -2515 -11788 -2279 -11787
<< metal5 >>
rect -3908 -3116 -3540 -3092
rect -3908 -3436 -3884 -3116
rect -3564 -3436 -3540 -3116
rect -3908 -3460 -3540 -3436
rect -3884 -4310 -3564 -3460
rect -2954 -4204 -2586 -4180
rect -2954 -4310 -2930 -4204
rect -3884 -4334 -2930 -4310
rect -2610 -4310 -2586 -4204
rect -3884 -4606 -2946 -4334
rect -2610 -4524 -2476 -4310
rect -2674 -4606 -2476 -4524
rect -3884 -4630 -2476 -4606
rect -2795 -6454 -2476 -4630
rect -2848 -6478 -2476 -6454
rect -2848 -6798 -2824 -6478
rect -2504 -6798 -2476 -6478
rect -2848 -6822 -2476 -6798
rect -2795 -10038 -2476 -6822
rect -3343 -10357 -2476 -10038
rect -3343 -14868 -3024 -10357
rect -2539 -11552 -2255 -11528
rect -2539 -11788 -2515 -11552
rect -2279 -11788 -2255 -11552
rect -2539 -11812 -2255 -11788
rect -2478 -12586 -2317 -11812
rect -3343 -15187 -2483 -14868
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -15016 0 1 -5376
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_1
timestamp 1695852000
transform 1 0 -17016 0 1 -5376
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_2
timestamp 1695852000
transform 1 0 19484 0 1 -5576
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_3
timestamp 1695852000
transform 1 0 17484 0 1 -5576
box -184 -124 1528 1016
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -4436 0 1 -6216
box -184 -124 1528 1592
use CNRATR_NCH_8C4F0  CNRATR_NCH_8C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -17016 0 1 -6776
box -184 -124 1912 1016
use CNRATR_NCH_8C4F0  CNRATR_NCH_8C4F0_1
timestamp 1695852000
transform 1 0 17484 0 1 -6976
box -184 -124 1912 1016
use CNRATR_NCH_8C12F0  CNRATR_NCH_8C12F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -17036 0 1 -9476
box -184 -124 1912 2168
use CNRATR_NCH_8C12F0  CNRATR_NCH_8C12F0_1
timestamp 1695852000
transform 1 0 17484 0 1 -9676
box -184 -124 1912 2168
use CNRATR_PCH_2C12F0  CNRATR_PCH_2C12F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -4316 0 1 -4296
box -184 -124 1336 2168
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 -11016 0 1 -3176
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_1
timestamp 1695852000
transform 1 0 -13016 0 1 -3176
box -184 -124 1528 1016
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 19484 0 1 -3876
box -184 -124 1528 1592
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_1
timestamp 1695852000
transform 1 0 17484 0 1 -3878
box -184 -124 1528 1592
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_2
timestamp 1695852000
transform 1 0 -17016 0 1 -3678
box -184 -124 1528 1592
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_3
timestamp 1695852000
transform 1 0 -15016 0 1 -3676
box -184 -124 1528 1592
use sky130_fd_pr__cap_mim_m3_2_BESJ5K  sky130_fd_pr__cap_mim_m3_2_BESJ5K_0
timestamp 1713440215
transform 0 -1 4122 1 0 -14771
box -2349 -6600 2371 6600
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 1 1288 0 1 1288
timestamp 1705271942
transform 1 0 -14660 0 1 -10700
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
array 0 3 1288 0 1 1288
timestamp 1705271942
transform 1 0 -10500 0 1 -10700
box 0 0 1340 1340
use SUNTR_RPPO2  SUNTR_RPPO2_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1713272488
transform 1 0 -13200 0 1 -7800
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_1
timestamp 1713272488
transform 1 0 -7600 0 1 -7800
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_2
timestamp 1713272488
transform 1 0 -10400 0 1 -7800
box 0 0 2672 4236
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712309819
transform 0 -1 17064 1 0 -10844
box 0 0 8720 4236
use SUNTR_RPPO16  SUNTR_RPPO16_1
timestamp 1712309819
transform 0 -1 1936 1 0 -10800
box 0 0 8720 4236
use SUNTR_RPPO16  SUNTR_RPPO16_2
timestamp 1712309819
transform 0 -1 -17436 1 0 -10644
box 0 0 8720 4236
use SUNTR_RPPO16  SUNTR_RPPO16_3
timestamp 1712309819
transform 0 -1 11236 1 0 -10800
box 0 0 8720 4236
use SUNTR_RPPO16  SUNTR_RPPO16_4
timestamp 1712309819
transform 0 -1 6736 1 0 -10800
box 0 0 8720 4236
<< labels >>
flabel metal1 -19760 -1540 16740 -1240 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel locali -21792 -11810 -3712 -11218 0 FreeSans 1600 0 0 0 VSS
port 6 nsew
flabel metal1 -2512 -4530 -2448 -2806 0 FreeSans 1600 0 0 0 RESET
port 3 nsew
flabel metal1 20060 -4750 20124 -3178 0 FreeSans 1600 0 0 0 COMPERATOR
port 25 nsew
<< end >>

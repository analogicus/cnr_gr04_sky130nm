magic
tech sky130B
magscale 1 2
timestamp 1713440215
<< error_p >>
rect -1951 160 -1583 184
rect -453 160 -85 184
rect 1045 160 1413 184
rect -1951 -160 -1927 160
rect -453 -160 -429 160
rect 1045 -160 1069 160
rect -1951 -184 -1583 -160
rect -453 -184 -85 -160
rect 1045 -184 1413 -160
<< metal4 >>
rect -2047 239 -949 280
rect -2047 -239 -1205 239
rect -969 -239 -949 239
rect -2047 -280 -949 -239
rect -549 239 549 280
rect -549 -239 293 239
rect 529 -239 549 239
rect -549 -280 549 -239
rect 949 239 2047 280
rect 949 -239 1791 239
rect 2027 -239 2047 239
rect 949 -280 2047 -239
<< via4 >>
rect -1205 -239 -969 239
rect 293 -239 529 239
rect 1791 -239 2027 239
<< mimcap2 >>
rect -1967 160 -1567 200
rect -1967 -160 -1927 160
rect -1607 -160 -1567 160
rect -1967 -200 -1567 -160
rect -469 160 -69 200
rect -469 -160 -429 160
rect -109 -160 -69 160
rect -469 -200 -69 -160
rect 1029 160 1429 200
rect 1029 -160 1069 160
rect 1389 -160 1429 160
rect 1029 -200 1429 -160
<< mimcap2contact >>
rect -1927 -160 -1607 160
rect -429 -160 -109 160
rect 1069 -160 1389 160
<< metal5 >>
rect -1247 239 -927 281
rect -1951 160 -1583 184
rect -1951 -160 -1927 160
rect -1607 -160 -1583 160
rect -1951 -184 -1583 -160
rect -1247 -239 -1205 239
rect -969 -239 -927 239
rect 251 239 571 281
rect -453 160 -85 184
rect -453 -160 -429 160
rect -109 -160 -85 160
rect -453 -184 -85 -160
rect -1247 -281 -927 -239
rect 251 -239 293 239
rect 529 -239 571 239
rect 1749 239 2069 281
rect 1045 160 1413 184
rect 1045 -160 1069 160
rect 1389 -160 1413 160
rect 1045 -184 1413 -160
rect 251 -281 571 -239
rect 1749 -239 1791 239
rect 2027 -239 2069 239
rect 1749 -281 2069 -239
<< properties >>
string FIXED_BBOX 949 -280 1509 280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

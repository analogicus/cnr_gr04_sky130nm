magic
tech sky130B
magscale 1 2
timestamp 1713460579
<< metal4 >>
rect -2349 6439 2349 6480
rect -2349 2361 2093 6439
rect 2329 2361 2349 6439
rect -2349 2320 2349 2361
rect -2349 2039 2349 2080
rect -2349 -2039 2093 2039
rect 2329 -2039 2349 2039
rect -2349 -2080 2349 -2039
rect -2349 -2361 2349 -2320
rect -2349 -6439 2093 -2361
rect 2329 -6439 2349 -2361
rect -2349 -6480 2349 -6439
<< via4 >>
rect 2093 2361 2329 6439
rect 2093 -2039 2329 2039
rect 2093 -6439 2329 -2361
<< mimcap2 >>
rect -2269 6360 1731 6400
rect -2269 2440 -2229 6360
rect 1691 2440 1731 6360
rect -2269 2400 1731 2440
rect -2269 1960 1731 2000
rect -2269 -1960 -2229 1960
rect 1691 -1960 1731 1960
rect -2269 -2000 1731 -1960
rect -2269 -2440 1731 -2400
rect -2269 -6360 -2229 -2440
rect 1691 -6360 1731 -2440
rect -2269 -6400 1731 -6360
<< mimcap2contact >>
rect -2229 2440 1691 6360
rect -2229 -1960 1691 1960
rect -2229 -6360 1691 -2440
<< metal5 >>
rect -429 6384 -109 6600
rect 2051 6439 2371 6600
rect -2253 6360 1715 6384
rect -2253 2440 -2229 6360
rect 1691 2440 1715 6360
rect -2253 2416 1715 2440
rect -429 1984 -109 2416
rect 2051 2361 2093 6439
rect 2329 2361 2371 6439
rect 2051 2039 2371 2361
rect -2253 1960 1715 1984
rect -2253 -1960 -2229 1960
rect 1691 -1960 1715 1960
rect -2253 -1984 1715 -1960
rect -429 -2416 -109 -1984
rect 2051 -2039 2093 2039
rect 2329 -2039 2371 2039
rect 2051 -2361 2371 -2039
rect -2253 -2440 1715 -2416
rect -2253 -6360 -2229 -2440
rect 1691 -6360 1715 -2440
rect -2253 -6384 1715 -6360
rect -429 -6600 -109 -6384
rect 2051 -6439 2093 -2361
rect 2329 -6439 2371 -2361
rect 2051 -6600 2371 -6439
<< properties >>
string FIXED_BBOX -2349 2320 1811 6480
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20.00 l 20.00 val 815.2 carea 2.00 cperi 0.19 nx 1 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1712916783
<< viali >>
rect 7573 9605 7607 9639
rect 7205 9537 7239 9571
rect 7021 9469 7055 9503
rect 6377 9333 6411 9367
rect 3525 8925 3559 8959
rect 4445 8925 4479 8959
rect 5917 8925 5951 8959
rect 7297 8925 7331 8959
rect 3280 8857 3314 8891
rect 4712 8857 4746 8891
rect 2145 8789 2179 8823
rect 5825 8789 5859 8823
rect 6561 8789 6595 8823
rect 6653 8789 6687 8823
rect 3893 8585 3927 8619
rect 5733 8585 5767 8619
rect 3617 8517 3651 8551
rect 1409 8449 1443 8483
rect 1676 8449 1710 8483
rect 3065 8449 3099 8483
rect 3249 8449 3283 8483
rect 3341 8449 3375 8483
rect 3525 8449 3559 8483
rect 3709 8449 3743 8483
rect 4445 8449 4479 8483
rect 6377 8449 6411 8483
rect 6644 8449 6678 8483
rect 2789 8313 2823 8347
rect 2973 8245 3007 8279
rect 7757 8245 7791 8279
rect 1593 8041 1627 8075
rect 2697 8041 2731 8075
rect 3065 8041 3099 8075
rect 4077 8041 4111 8075
rect 4445 8041 4479 8075
rect 6929 8041 6963 8075
rect 3157 7973 3191 8007
rect 5825 7905 5859 7939
rect 6285 7905 6319 7939
rect 1777 7837 1811 7871
rect 1961 7837 1995 7871
rect 2605 7837 2639 7871
rect 2881 7837 2915 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 3617 7837 3651 7871
rect 3893 7837 3927 7871
rect 4353 7837 4387 7871
rect 5089 7837 5123 7871
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 5457 7837 5491 7871
rect 5549 7837 5583 7871
rect 8309 7837 8343 7871
rect 4261 7769 4295 7803
rect 3525 7701 3559 7735
rect 8493 7701 8527 7735
rect 1869 7497 1903 7531
rect 5549 7497 5583 7531
rect 6469 7497 6503 7531
rect 1501 7429 1535 7463
rect 1685 7429 1719 7463
rect 3868 7429 3902 7463
rect 4077 7429 4111 7463
rect 2237 7361 2271 7395
rect 2973 7361 3007 7395
rect 3617 7361 3651 7395
rect 4353 7361 4387 7395
rect 4445 7361 4479 7395
rect 6193 7361 6227 7395
rect 6561 7361 6595 7395
rect 7021 7361 7055 7395
rect 7277 7361 7311 7395
rect 2329 7293 2363 7327
rect 2513 7293 2547 7327
rect 3985 7293 4019 7327
rect 4721 7293 4755 7327
rect 4905 7293 4939 7327
rect 4629 7225 4663 7259
rect 3709 7157 3743 7191
rect 4537 7157 4571 7191
rect 5457 7157 5491 7191
rect 8401 7157 8435 7191
rect 2973 6953 3007 6987
rect 3157 6953 3191 6987
rect 4169 6953 4203 6987
rect 3249 6885 3283 6919
rect 1593 6817 1627 6851
rect 3617 6817 3651 6851
rect 6377 6817 6411 6851
rect 7205 6817 7239 6851
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 5917 6749 5951 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 6561 6749 6595 6783
rect 7021 6749 7055 6783
rect 7113 6749 7147 6783
rect 1860 6681 1894 6715
rect 5282 6681 5316 6715
rect 5733 6681 5767 6715
rect 6837 6681 6871 6715
rect 7450 6681 7484 6715
rect 6101 6613 6135 6647
rect 6745 6613 6779 6647
rect 6929 6613 6963 6647
rect 8585 6613 8619 6647
rect 1777 6409 1811 6443
rect 2697 6409 2731 6443
rect 5365 6409 5399 6443
rect 6577 6409 6611 6443
rect 7205 6409 7239 6443
rect 3700 6341 3734 6375
rect 6377 6341 6411 6375
rect 6837 6341 6871 6375
rect 7037 6341 7071 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2053 6273 2087 6307
rect 3433 6273 3467 6307
rect 4997 6273 5031 6307
rect 5181 6273 5215 6307
rect 8309 6273 8343 6307
rect 2789 6205 2823 6239
rect 2881 6205 2915 6239
rect 4905 6205 4939 6239
rect 2329 6137 2363 6171
rect 4813 6137 4847 6171
rect 8493 6137 8527 6171
rect 1501 6069 1535 6103
rect 6561 6069 6595 6103
rect 6745 6069 6779 6103
rect 7021 6069 7055 6103
rect 2605 5865 2639 5899
rect 2881 5865 2915 5899
rect 5641 5865 5675 5899
rect 6561 5865 6595 5899
rect 6837 5865 6871 5899
rect 3249 5797 3283 5831
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 1778 5661 1812 5695
rect 1961 5661 1995 5695
rect 2191 5661 2225 5695
rect 3065 5661 3099 5695
rect 3157 5661 3191 5695
rect 3893 5661 3927 5695
rect 4077 5661 4111 5695
rect 4353 5661 4387 5695
rect 6469 5661 6503 5695
rect 6561 5661 6595 5695
rect 7941 5661 7975 5695
rect 8309 5661 8343 5695
rect 2053 5593 2087 5627
rect 2421 5593 2455 5627
rect 6805 5593 6839 5627
rect 7021 5593 7055 5627
rect 1593 5525 1627 5559
rect 2329 5525 2363 5559
rect 2621 5525 2655 5559
rect 2789 5525 2823 5559
rect 3985 5525 4019 5559
rect 6193 5525 6227 5559
rect 6653 5525 6687 5559
rect 8125 5525 8159 5559
rect 8493 5525 8527 5559
rect 1501 5321 1535 5355
rect 2329 5321 2363 5355
rect 3801 5321 3835 5355
rect 5365 5321 5399 5355
rect 6193 5321 6227 5355
rect 6929 5321 6963 5355
rect 8493 5321 8527 5355
rect 2688 5253 2722 5287
rect 5641 5253 5675 5287
rect 5825 5253 5859 5287
rect 6041 5253 6075 5287
rect 6377 5253 6411 5287
rect 6561 5253 6595 5287
rect 7358 5253 7392 5287
rect 1593 5185 1627 5219
rect 1685 5185 1719 5219
rect 4077 5185 4111 5219
rect 5089 5185 5123 5219
rect 5365 5185 5399 5219
rect 6745 5185 6779 5219
rect 6837 5185 6871 5219
rect 7021 5185 7055 5219
rect 2421 5117 2455 5151
rect 4721 5117 4755 5151
rect 4813 5117 4847 5151
rect 5457 5117 5491 5151
rect 7113 5117 7147 5151
rect 5273 5049 5307 5083
rect 4905 4981 4939 5015
rect 6009 4981 6043 5015
rect 1409 4777 1443 4811
rect 4629 4777 4663 4811
rect 4997 4777 5031 4811
rect 5641 4777 5675 4811
rect 8585 4777 8619 4811
rect 5089 4709 5123 4743
rect 4353 4641 4387 4675
rect 7205 4641 7239 4675
rect 2522 4573 2556 4607
rect 2789 4573 2823 4607
rect 4169 4573 4203 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 4721 4573 4755 4607
rect 4905 4573 4939 4607
rect 5181 4573 5215 4607
rect 5549 4573 5583 4607
rect 5733 4573 5767 4607
rect 6469 4573 6503 4607
rect 6653 4573 6687 4607
rect 6745 4573 6779 4607
rect 6837 4573 6871 4607
rect 7113 4505 7147 4539
rect 7450 4505 7484 4539
rect 5457 4437 5491 4471
rect 4997 4233 5031 4267
rect 6561 4233 6595 4267
rect 4537 4165 4571 4199
rect 5365 4165 5399 4199
rect 3157 4097 3191 4131
rect 3341 4097 3375 4131
rect 3433 4097 3467 4131
rect 4997 4097 5031 4131
rect 5181 4097 5215 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 8493 4097 8527 4131
rect 6745 4029 6779 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7849 4029 7883 4063
rect 4353 3961 4387 3995
rect 4905 3961 4939 3995
rect 3157 3893 3191 3927
rect 4537 3893 4571 3927
rect 7297 3893 7331 3927
rect 3985 3689 4019 3723
rect 3893 3621 3927 3655
rect 8493 3621 8527 3655
rect 3525 3553 3559 3587
rect 4077 3553 4111 3587
rect 6101 3553 6135 3587
rect 3801 3485 3835 3519
rect 4353 3485 4387 3519
rect 8309 3485 8343 3519
rect 2973 3349 3007 3383
rect 4353 3145 4387 3179
rect 4712 3077 4746 3111
rect 5917 3077 5951 3111
rect 6377 3077 6411 3111
rect 6577 3077 6611 3111
rect 2329 3009 2363 3043
rect 2596 3009 2630 3043
rect 4445 3009 4479 3043
rect 6101 3009 6135 3043
rect 6193 3009 6227 3043
rect 6837 3009 6871 3043
rect 7093 3009 7127 3043
rect 3893 2941 3927 2975
rect 3985 2941 4019 2975
rect 4077 2941 4111 2975
rect 4169 2941 4203 2975
rect 6745 2873 6779 2907
rect 3709 2805 3743 2839
rect 5825 2805 5859 2839
rect 6193 2805 6227 2839
rect 6561 2805 6595 2839
rect 8217 2805 8251 2839
rect 1501 2601 1535 2635
rect 5089 2601 5123 2635
rect 5733 2601 5767 2635
rect 6377 2601 6411 2635
rect 4445 2465 4479 2499
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 3617 2397 3651 2431
rect 3893 2397 3927 2431
rect 4537 2397 4571 2431
rect 5549 2397 5583 2431
rect 5641 2397 5675 2431
rect 6561 2397 6595 2431
rect 6837 2397 6871 2431
rect 2636 2329 2670 2363
rect 4721 2329 4755 2363
rect 3065 2261 3099 2295
rect 3433 2261 3467 2295
rect 4813 2261 4847 2295
rect 4905 2261 4939 2295
rect 5365 2261 5399 2295
rect 6745 2261 6779 2295
<< metal1 >>
rect 1104 9818 8924 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 8924 9818
rect 1104 9744 8924 9766
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 7561 9639 7619 9645
rect 7561 9636 7573 9639
rect 5868 9608 7573 9636
rect 5868 9596 5874 9608
rect 7561 9605 7573 9608
rect 7607 9605 7619 9639
rect 7561 9599 7619 9605
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 6236 9540 7205 9568
rect 6236 9528 6242 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9500 7067 9503
rect 7282 9500 7288 9512
rect 7055 9472 7288 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 6362 9324 6368 9376
rect 6420 9324 6426 9376
rect 1104 9274 8924 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 8924 9274
rect 1104 9200 8924 9222
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 2188 8928 3525 8956
rect 2188 8916 2194 8928
rect 3513 8925 3525 8928
rect 3559 8956 3571 8959
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 3559 8928 4445 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 4433 8925 4445 8928
rect 4479 8956 4491 8959
rect 5718 8956 5724 8968
rect 4479 8928 5724 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 5905 8959 5963 8965
rect 5905 8956 5917 8959
rect 5828 8928 5917 8956
rect 3268 8891 3326 8897
rect 3268 8857 3280 8891
rect 3314 8888 3326 8891
rect 3878 8888 3884 8900
rect 3314 8860 3884 8888
rect 3314 8857 3326 8860
rect 3268 8851 3326 8857
rect 3878 8848 3884 8860
rect 3936 8848 3942 8900
rect 4706 8897 4712 8900
rect 4700 8851 4712 8897
rect 4706 8848 4712 8851
rect 4764 8848 4770 8900
rect 2133 8823 2191 8829
rect 2133 8789 2145 8823
rect 2179 8820 2191 8823
rect 2590 8820 2596 8832
rect 2179 8792 2596 8820
rect 2179 8789 2191 8792
rect 2133 8783 2191 8789
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 5828 8829 5856 8928
rect 5905 8925 5917 8928
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5316 8792 5825 8820
rect 5316 8780 5322 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 5960 8792 6561 8820
rect 5960 8780 5966 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 6638 8780 6644 8832
rect 6696 8780 6702 8832
rect 1104 8730 8924 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8924 8730
rect 1104 8656 8924 8678
rect 2130 8576 2136 8628
rect 2188 8576 2194 8628
rect 3878 8576 3884 8628
rect 3936 8576 3942 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 2148 8548 2176 8576
rect 1412 8520 2176 8548
rect 3605 8551 3663 8557
rect 1412 8492 1440 8520
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 5534 8548 5540 8560
rect 3651 8520 5540 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1670 8489 1676 8492
rect 1664 8443 1676 8489
rect 1670 8440 1676 8443
rect 1728 8440 1734 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3068 8344 3096 8443
rect 3142 8440 3148 8492
rect 3200 8440 3206 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8449 3387 8483
rect 3329 8443 3387 8449
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 5626 8480 5632 8492
rect 4479 8452 5632 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 3160 8412 3188 8440
rect 3344 8412 3372 8443
rect 3160 8384 3372 8412
rect 2823 8316 3096 8344
rect 3528 8344 3556 8443
rect 3712 8412 3740 8443
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5736 8480 5764 8576
rect 6914 8548 6920 8560
rect 6380 8520 6920 8548
rect 6380 8489 6408 8520
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 5736 8452 6377 8480
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6632 8483 6690 8489
rect 6632 8449 6644 8483
rect 6678 8480 6690 8483
rect 7006 8480 7012 8492
rect 6678 8452 7012 8480
rect 6678 8449 6690 8452
rect 6632 8443 6690 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 4614 8412 4620 8424
rect 3712 8384 4620 8412
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 5902 8344 5908 8356
rect 3528 8316 5908 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 2792 8276 2820 8307
rect 2372 8248 2820 8276
rect 2372 8236 2378 8248
rect 2958 8236 2964 8288
rect 3016 8236 3022 8288
rect 3068 8276 3096 8316
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 4062 8276 4068 8288
rect 3068 8248 4068 8276
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 7282 8276 7288 8288
rect 4948 8248 7288 8276
rect 4948 8236 4954 8248
rect 7282 8236 7288 8248
rect 7340 8276 7346 8288
rect 7745 8279 7803 8285
rect 7745 8276 7757 8279
rect 7340 8248 7757 8276
rect 7340 8236 7346 8248
rect 7745 8245 7757 8248
rect 7791 8245 7803 8279
rect 7745 8239 7803 8245
rect 1104 8186 8924 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 8924 8186
rect 1104 8112 8924 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1670 8072 1676 8084
rect 1627 8044 1676 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 2958 8072 2964 8084
rect 2731 8044 2964 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3234 8072 3240 8084
rect 3099 8044 3240 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3234 8032 3240 8044
rect 3292 8032 3298 8084
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 4246 8072 4252 8084
rect 4111 8044 4252 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4614 8072 4620 8084
rect 4479 8044 4620 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 4706 8032 4712 8084
rect 4764 8032 4770 8084
rect 5166 8072 5172 8084
rect 4816 8044 5172 8072
rect 2590 7964 2596 8016
rect 2648 8004 2654 8016
rect 3145 8007 3203 8013
rect 2648 7976 2774 8004
rect 2648 7964 2654 7976
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 2038 7868 2044 7880
rect 1995 7840 2044 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2590 7828 2596 7880
rect 2648 7828 2654 7880
rect 2746 7868 2774 7976
rect 3145 7973 3157 8007
rect 3191 8004 3203 8007
rect 4724 8004 4752 8032
rect 3191 7976 4752 8004
rect 3191 7973 3203 7976
rect 3145 7967 3203 7973
rect 4522 7936 4528 7948
rect 3620 7908 4528 7936
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2746 7840 2881 7868
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3050 7828 3056 7880
rect 3108 7868 3114 7880
rect 3620 7877 3648 7908
rect 4522 7896 4528 7908
rect 4580 7936 4586 7948
rect 4816 7936 4844 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7006 8072 7012 8084
rect 6963 8044 7012 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 5258 7936 5264 7948
rect 4580 7908 4844 7936
rect 5000 7908 5264 7936
rect 4580 7896 4586 7908
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 3108 7840 3249 7868
rect 3108 7828 3114 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3881 7871 3939 7877
rect 3881 7837 3893 7871
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4706 7868 4712 7880
rect 4387 7840 4712 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 3344 7800 3372 7831
rect 3200 7772 3372 7800
rect 3200 7760 3206 7772
rect 3510 7692 3516 7744
rect 3568 7692 3574 7744
rect 3896 7732 3924 7831
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4249 7803 4307 7809
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 5000 7800 5028 7908
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 5718 7936 5724 7948
rect 5368 7908 5724 7936
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 4295 7772 5028 7800
rect 5092 7800 5120 7831
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5368 7877 5396 7908
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7936 5871 7939
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 5859 7908 6285 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 5534 7828 5540 7880
rect 5592 7868 5598 7880
rect 6362 7868 6368 7880
rect 5592 7840 6368 7868
rect 5592 7828 5598 7840
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7064 7840 8309 7868
rect 7064 7828 7070 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 6178 7800 6184 7812
rect 5092 7772 6184 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 3970 7732 3976 7744
rect 3896 7704 3976 7732
rect 3970 7692 3976 7704
rect 4028 7732 4034 7744
rect 5092 7732 5120 7772
rect 6178 7760 6184 7772
rect 6236 7760 6242 7812
rect 4028 7704 5120 7732
rect 4028 7692 4034 7704
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 1104 7642 8924 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8924 7642
rect 1104 7568 8924 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 1857 7531 1915 7537
rect 1857 7528 1869 7531
rect 1820 7500 1869 7528
rect 1820 7488 1826 7500
rect 1857 7497 1869 7500
rect 1903 7497 1915 7531
rect 1857 7491 1915 7497
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2096 7500 3464 7528
rect 2096 7488 2102 7500
rect 1210 7420 1216 7472
rect 1268 7460 1274 7472
rect 1489 7463 1547 7469
rect 1489 7460 1501 7463
rect 1268 7432 1501 7460
rect 1268 7420 1274 7432
rect 1489 7429 1501 7432
rect 1535 7429 1547 7463
rect 1489 7423 1547 7429
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 2774 7460 2780 7472
rect 1719 7432 2780 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 2774 7420 2780 7432
rect 2832 7460 2838 7472
rect 3050 7460 3056 7472
rect 2832 7432 3056 7460
rect 2832 7420 2838 7432
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 3436 7460 3464 7500
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 3568 7500 5028 7528
rect 3568 7488 3574 7500
rect 3856 7463 3914 7469
rect 3856 7460 3868 7463
rect 3436 7432 3868 7460
rect 3856 7429 3868 7432
rect 3902 7429 3914 7463
rect 3856 7423 3914 7429
rect 4062 7420 4068 7472
rect 4120 7420 4126 7472
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 4706 7460 4712 7472
rect 4304 7432 4712 7460
rect 4304 7420 4310 7432
rect 2222 7352 2228 7404
rect 2280 7352 2286 7404
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 4448 7401 4476 7432
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 5000 7460 5028 7500
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5500 7500 5549 7528
rect 5500 7488 5506 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5537 7491 5595 7497
rect 5644 7500 6469 7528
rect 5644 7460 5672 7500
rect 6457 7497 6469 7500
rect 6503 7497 6515 7531
rect 6457 7491 6515 7497
rect 5000 7432 5672 7460
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2648 7364 2973 7392
rect 2648 7352 2654 7364
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7392 3663 7395
rect 4341 7395 4399 7401
rect 4341 7392 4353 7395
rect 3651 7364 4353 7392
rect 3651 7361 3663 7364
rect 3605 7355 3663 7361
rect 4341 7361 4353 7364
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 1946 7284 1952 7336
rect 2004 7324 2010 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 2004 7296 2329 7324
rect 2004 7284 2010 7296
rect 2317 7293 2329 7296
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7324 2559 7327
rect 2682 7324 2688 7336
rect 2547 7296 2688 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 2682 7284 2688 7296
rect 2740 7324 2746 7336
rect 3973 7327 4031 7333
rect 2740 7284 2774 7324
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 2746 7256 2774 7284
rect 3988 7256 4016 7287
rect 2746 7228 4016 7256
rect 4540 7256 4568 7352
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7293 4767 7327
rect 4709 7287 4767 7293
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5350 7324 5356 7336
rect 4939 7296 5356 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 4617 7259 4675 7265
rect 4617 7256 4629 7259
rect 4540 7228 4629 7256
rect 4617 7225 4629 7228
rect 4663 7225 4675 7259
rect 4724 7256 4752 7287
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5920 7324 5948 7352
rect 6564 7324 6592 7355
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6972 7364 7021 7392
rect 6972 7352 6978 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 5920 7296 6592 7324
rect 6638 7284 6644 7336
rect 6696 7284 6702 7336
rect 6656 7256 6684 7284
rect 4724 7228 6684 7256
rect 4617 7219 4675 7225
rect 3694 7148 3700 7200
rect 3752 7148 3758 7200
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 3844 7160 4537 7188
rect 3844 7148 3850 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4525 7151 4583 7157
rect 5442 7148 5448 7200
rect 5500 7148 5506 7200
rect 7024 7188 7052 7355
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7265 7395 7323 7401
rect 7265 7392 7277 7395
rect 7156 7364 7277 7392
rect 7156 7352 7162 7364
rect 7265 7361 7277 7364
rect 7311 7361 7323 7395
rect 7265 7355 7323 7361
rect 7190 7188 7196 7200
rect 7024 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 1104 7098 8924 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 8924 7098
rect 1104 7024 8924 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 2961 6987 3019 6993
rect 2961 6984 2973 6987
rect 2648 6956 2973 6984
rect 2648 6944 2654 6956
rect 2961 6953 2973 6956
rect 3007 6953 3019 6987
rect 2961 6947 3019 6953
rect 3142 6944 3148 6996
rect 3200 6984 3206 6996
rect 3786 6984 3792 6996
rect 3200 6956 3792 6984
rect 3200 6944 3206 6956
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4157 6987 4215 6993
rect 4157 6984 4169 6987
rect 4028 6956 4169 6984
rect 4028 6944 4034 6956
rect 4157 6953 4169 6956
rect 4203 6953 4215 6987
rect 4157 6947 4215 6953
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 3237 6919 3295 6925
rect 3237 6916 3249 6919
rect 2740 6888 3249 6916
rect 2740 6876 2746 6888
rect 3237 6885 3249 6888
rect 3283 6885 3295 6919
rect 3237 6879 3295 6885
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1581 6851 1639 6857
rect 1581 6848 1593 6851
rect 1452 6820 1593 6848
rect 1452 6808 1458 6820
rect 1581 6817 1593 6820
rect 1627 6817 1639 6851
rect 1581 6811 1639 6817
rect 3605 6851 3663 6857
rect 3605 6817 3617 6851
rect 3651 6848 3663 6851
rect 3988 6848 4016 6944
rect 6454 6876 6460 6928
rect 6512 6916 6518 6928
rect 7006 6916 7012 6928
rect 6512 6888 7012 6916
rect 6512 6876 6518 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 3651 6820 4016 6848
rect 5920 6820 6377 6848
rect 3651 6817 3663 6820
rect 3605 6811 3663 6817
rect 1596 6780 1624 6811
rect 3418 6780 3424 6792
rect 1596 6752 3424 6780
rect 3418 6740 3424 6752
rect 3476 6780 3482 6792
rect 5920 6789 5948 6820
rect 6365 6817 6377 6820
rect 6411 6848 6423 6851
rect 6411 6820 7144 6848
rect 6411 6817 6423 6820
rect 6365 6811 6423 6817
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 3476 6752 5549 6780
rect 3476 6740 3482 6752
rect 5537 6749 5549 6752
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 1854 6721 1860 6724
rect 1848 6675 1860 6721
rect 1854 6672 1860 6675
rect 1912 6672 1918 6724
rect 5258 6672 5264 6724
rect 5316 6721 5322 6724
rect 5316 6675 5328 6721
rect 5644 6712 5672 6743
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 5552 6684 5672 6712
rect 5721 6715 5779 6721
rect 5316 6672 5322 6675
rect 5552 6656 5580 6684
rect 5721 6681 5733 6715
rect 5767 6712 5779 6715
rect 6472 6712 6500 6740
rect 5767 6684 6500 6712
rect 6564 6712 6592 6743
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6696 6752 6960 6780
rect 6696 6740 6702 6752
rect 6822 6712 6828 6724
rect 6564 6684 6828 6712
rect 5767 6681 5779 6684
rect 5721 6675 5779 6681
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 5534 6604 5540 6656
rect 5592 6604 5598 6656
rect 6086 6604 6092 6656
rect 6144 6604 6150 6656
rect 6730 6604 6736 6656
rect 6788 6604 6794 6656
rect 6932 6653 6960 6752
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7116 6789 7144 6820
rect 7190 6808 7196 6860
rect 7248 6808 7254 6860
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6780 7159 6783
rect 7282 6780 7288 6792
rect 7147 6752 7288 6780
rect 7147 6749 7159 6752
rect 7101 6743 7159 6749
rect 7282 6740 7288 6752
rect 7340 6780 7346 6792
rect 8386 6780 8392 6792
rect 7340 6752 8392 6780
rect 7340 6740 7346 6752
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7438 6715 7496 6721
rect 7438 6712 7450 6715
rect 7248 6684 7450 6712
rect 7248 6672 7254 6684
rect 7438 6681 7450 6684
rect 7484 6681 7496 6715
rect 7438 6675 7496 6681
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 8570 6604 8576 6656
rect 8628 6604 8634 6656
rect 1104 6554 8924 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8924 6554
rect 1104 6480 8924 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 1854 6440 1860 6452
rect 1811 6412 1860 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 2590 6400 2596 6452
rect 2648 6440 2654 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2648 6412 2697 6440
rect 2648 6400 2654 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 3418 6400 3424 6452
rect 3476 6400 3482 6452
rect 5258 6400 5264 6452
rect 5316 6440 5322 6452
rect 5353 6443 5411 6449
rect 5353 6440 5365 6443
rect 5316 6412 5365 6440
rect 5316 6400 5322 6412
rect 5353 6409 5365 6412
rect 5399 6409 5411 6443
rect 5353 6403 5411 6409
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 6565 6443 6623 6449
rect 6565 6440 6577 6443
rect 6144 6412 6577 6440
rect 6144 6400 6150 6412
rect 6565 6409 6577 6412
rect 6611 6409 6623 6443
rect 6565 6403 6623 6409
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 6788 6412 7144 6440
rect 6788 6400 6794 6412
rect 1670 6264 1676 6316
rect 1728 6264 1734 6316
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1964 6168 1992 6267
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 3436 6313 3464 6400
rect 3694 6381 3700 6384
rect 3688 6372 3700 6381
rect 3655 6344 3700 6372
rect 3688 6335 3700 6344
rect 3694 6332 3700 6335
rect 3752 6332 3758 6384
rect 5718 6372 5724 6384
rect 5184 6344 5724 6372
rect 3421 6307 3479 6313
rect 2740 6276 2912 6304
rect 2740 6264 2746 6276
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 2884 6245 2912 6276
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4764 6276 4997 6304
rect 4764 6264 4770 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5184 6313 5212 6344
rect 5718 6332 5724 6344
rect 5776 6332 5782 6384
rect 6365 6375 6423 6381
rect 6365 6341 6377 6375
rect 6411 6372 6423 6375
rect 6825 6375 6883 6381
rect 6825 6372 6837 6375
rect 6411 6344 6837 6372
rect 6411 6341 6423 6344
rect 6365 6335 6423 6341
rect 6825 6341 6837 6344
rect 6871 6341 6883 6375
rect 6825 6335 6883 6341
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 5132 6276 5181 6304
rect 5132 6264 5138 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2280 6208 2789 6236
rect 2280 6196 2286 6208
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6236 4951 6239
rect 5460 6236 5488 6264
rect 4939 6208 5488 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 2317 6171 2375 6177
rect 2317 6168 2329 6171
rect 1964 6140 2329 6168
rect 2317 6137 2329 6140
rect 2363 6137 2375 6171
rect 2317 6131 2375 6137
rect 4801 6171 4859 6177
rect 4801 6137 4813 6171
rect 4847 6168 4859 6171
rect 5350 6168 5356 6180
rect 4847 6140 5356 6168
rect 4847 6137 4859 6140
rect 4801 6131 4859 6137
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 1486 6060 1492 6112
rect 1544 6060 1550 6112
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 2774 6100 2780 6112
rect 1912 6072 2780 6100
rect 1912 6060 1918 6072
rect 2774 6060 2780 6072
rect 2832 6100 2838 6112
rect 3142 6100 3148 6112
rect 2832 6072 3148 6100
rect 2832 6060 2838 6072
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 6380 6100 6408 6335
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 7025 6375 7083 6381
rect 7025 6372 7037 6375
rect 6972 6344 7037 6372
rect 6972 6332 6978 6344
rect 7025 6341 7037 6344
rect 7071 6341 7083 6375
rect 7025 6335 7083 6341
rect 7116 6304 7144 6412
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 8297 6307 8355 6313
rect 7116 6276 7236 6304
rect 6638 6196 6644 6248
rect 6696 6196 6702 6248
rect 7098 6236 7104 6248
rect 6932 6208 7104 6236
rect 4764 6072 6408 6100
rect 6549 6103 6607 6109
rect 4764 6060 4770 6072
rect 6549 6069 6561 6103
rect 6595 6100 6607 6103
rect 6656 6100 6684 6196
rect 6595 6072 6684 6100
rect 6733 6103 6791 6109
rect 6595 6069 6607 6072
rect 6549 6063 6607 6069
rect 6733 6069 6745 6103
rect 6779 6100 6791 6103
rect 6932 6100 6960 6208
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 6779 6072 6960 6100
rect 7009 6103 7067 6109
rect 6779 6069 6791 6072
rect 6733 6063 6791 6069
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7208 6100 7236 6276
rect 8297 6273 8309 6307
rect 8343 6304 8355 6307
rect 8386 6304 8392 6316
rect 8343 6276 8392 6304
rect 8343 6273 8355 6276
rect 8297 6267 8355 6273
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 8478 6128 8484 6180
rect 8536 6128 8542 6180
rect 7055 6072 7236 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 1104 6010 8924 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 8924 6010
rect 1104 5936 8924 5958
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 1636 5868 2605 5896
rect 1636 5856 1642 5868
rect 2593 5865 2605 5868
rect 2639 5896 2651 5899
rect 2869 5899 2927 5905
rect 2869 5896 2881 5899
rect 2639 5868 2881 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 2869 5865 2881 5868
rect 2915 5865 2927 5899
rect 2869 5859 2927 5865
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5626 5896 5632 5908
rect 4856 5868 5632 5896
rect 4856 5856 4862 5868
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6595 5868 6837 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6825 5865 6837 5868
rect 6871 5896 6883 5899
rect 7282 5896 7288 5908
rect 6871 5868 7288 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 8570 5856 8576 5908
rect 8628 5856 8634 5908
rect 2130 5788 2136 5840
rect 2188 5828 2194 5840
rect 3237 5831 3295 5837
rect 3237 5828 3249 5831
rect 2188 5800 3249 5828
rect 2188 5788 2194 5800
rect 3237 5797 3249 5800
rect 3283 5828 3295 5831
rect 5074 5828 5080 5840
rect 3283 5800 5080 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 1854 5760 1860 5772
rect 1688 5732 1860 5760
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1688 5701 1716 5732
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 1964 5732 5396 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1762 5652 1768 5704
rect 1820 5652 1826 5704
rect 1964 5701 1992 5732
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 2179 5695 2237 5701
rect 2179 5661 2191 5695
rect 2225 5692 2237 5695
rect 2314 5692 2320 5704
rect 2225 5664 2320 5692
rect 2225 5661 2237 5664
rect 2179 5655 2237 5661
rect 2314 5652 2320 5664
rect 2372 5652 2378 5704
rect 3050 5652 3056 5704
rect 3108 5652 3114 5704
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3881 5695 3939 5701
rect 3881 5692 3893 5695
rect 3200 5664 3893 5692
rect 3200 5652 3206 5664
rect 3881 5661 3893 5664
rect 3927 5661 3939 5695
rect 3881 5655 3939 5661
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4614 5692 4620 5704
rect 4387 5664 4620 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5368 5636 5396 5732
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 6328 5732 6960 5760
rect 6328 5720 6334 5732
rect 6472 5701 6500 5732
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 2038 5584 2044 5636
rect 2096 5584 2102 5636
rect 2409 5627 2467 5633
rect 2409 5624 2421 5627
rect 2148 5596 2421 5624
rect 2148 5568 2176 5596
rect 2409 5593 2421 5596
rect 2455 5593 2467 5627
rect 2409 5587 2467 5593
rect 5350 5584 5356 5636
rect 5408 5584 5414 5636
rect 6564 5624 6592 5652
rect 6793 5627 6851 5633
rect 6793 5624 6805 5627
rect 6564 5596 6805 5624
rect 6793 5593 6805 5596
rect 6839 5624 6851 5627
rect 6932 5624 6960 5732
rect 7300 5732 8340 5760
rect 7009 5627 7067 5633
rect 7009 5624 7021 5627
rect 6839 5593 6868 5624
rect 6932 5596 7021 5624
rect 6793 5587 6868 5593
rect 7009 5593 7021 5596
rect 7055 5624 7067 5627
rect 7300 5624 7328 5732
rect 8312 5701 8340 5732
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8588 5692 8616 5856
rect 8343 5664 8616 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 7055 5596 7328 5624
rect 7944 5624 7972 5655
rect 8570 5624 8576 5636
rect 7944 5596 8576 5624
rect 7055 5593 7067 5596
rect 7009 5587 7067 5593
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 1946 5556 1952 5568
rect 1627 5528 1952 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2130 5516 2136 5568
rect 2188 5516 2194 5568
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 2498 5556 2504 5568
rect 2363 5528 2504 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 2590 5516 2596 5568
rect 2648 5565 2654 5568
rect 2648 5559 2667 5565
rect 2655 5525 2667 5559
rect 2648 5519 2667 5525
rect 2648 5516 2654 5519
rect 2774 5516 2780 5568
rect 2832 5516 2838 5568
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 4706 5556 4712 5568
rect 4019 5528 4712 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 6181 5559 6239 5565
rect 6181 5556 6193 5559
rect 5684 5528 6193 5556
rect 5684 5516 5690 5528
rect 6181 5525 6193 5528
rect 6227 5525 6239 5559
rect 6181 5519 6239 5525
rect 6638 5516 6644 5568
rect 6696 5516 6702 5568
rect 6840 5556 6868 5587
rect 8570 5584 8576 5596
rect 8628 5584 8634 5636
rect 7098 5556 7104 5568
rect 6840 5528 7104 5556
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 8110 5516 8116 5568
rect 8168 5516 8174 5568
rect 8478 5516 8484 5568
rect 8536 5516 8542 5568
rect 1104 5466 8924 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8924 5466
rect 1104 5392 8924 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 2038 5352 2044 5364
rect 1535 5324 2044 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2590 5352 2596 5364
rect 2372 5324 2596 5352
rect 2372 5312 2378 5324
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 3789 5355 3847 5361
rect 3789 5321 3801 5355
rect 3835 5352 3847 5355
rect 3835 5324 4108 5352
rect 3835 5321 3847 5324
rect 3789 5315 3847 5321
rect 2676 5287 2734 5293
rect 2676 5253 2688 5287
rect 2722 5284 2734 5287
rect 2774 5284 2780 5296
rect 2722 5256 2780 5284
rect 2722 5253 2734 5256
rect 2676 5247 2734 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 4080 5228 4108 5324
rect 5350 5312 5356 5364
rect 5408 5312 5414 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6227 5324 6776 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 4706 5244 4712 5296
rect 4764 5284 4770 5296
rect 5166 5284 5172 5296
rect 4764 5256 5172 5284
rect 4764 5244 4770 5256
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5626 5244 5632 5296
rect 5684 5244 5690 5296
rect 5810 5244 5816 5296
rect 5868 5244 5874 5296
rect 6029 5287 6087 5293
rect 6029 5253 6041 5287
rect 6075 5284 6087 5287
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 6075 5256 6377 5284
rect 6075 5253 6087 5256
rect 6029 5247 6087 5253
rect 6365 5253 6377 5256
rect 6411 5253 6423 5287
rect 6365 5247 6423 5253
rect 6546 5244 6552 5296
rect 6604 5244 6610 5296
rect 6748 5284 6776 5324
rect 6914 5312 6920 5364
rect 6972 5312 6978 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 7156 5324 8493 5352
rect 7156 5312 7162 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 7346 5287 7404 5293
rect 7346 5284 7358 5287
rect 6748 5256 7358 5284
rect 7346 5253 7358 5256
rect 7392 5253 7404 5287
rect 7346 5247 7404 5253
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 1670 5176 1676 5228
rect 1728 5176 1734 5228
rect 4062 5176 4068 5228
rect 4120 5176 4126 5228
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5258 5216 5264 5228
rect 5123 5188 5264 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 5592 5188 6745 5216
rect 5592 5176 5598 5188
rect 6733 5185 6745 5188
rect 6779 5216 6791 5219
rect 6822 5216 6828 5228
rect 6779 5188 6828 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 2409 5111 2467 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4755 5120 4813 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 4801 5111 4859 5117
rect 2424 5012 2452 5111
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5040 5120 5457 5148
rect 5040 5108 5046 5120
rect 5445 5117 5457 5120
rect 5491 5148 5503 5151
rect 5902 5148 5908 5160
rect 5491 5120 5908 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 7024 5148 7052 5179
rect 6748 5120 7052 5148
rect 3510 5040 3516 5092
rect 3568 5080 3574 5092
rect 5261 5083 5319 5089
rect 5261 5080 5273 5083
rect 3568 5052 5273 5080
rect 3568 5040 3574 5052
rect 5261 5049 5273 5052
rect 5307 5049 5319 5083
rect 5261 5043 5319 5049
rect 6748 5024 6776 5120
rect 7098 5108 7104 5160
rect 7156 5108 7162 5160
rect 2774 5012 2780 5024
rect 2424 4984 2780 5012
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 4890 4972 4896 5024
rect 4948 4972 4954 5024
rect 5994 4972 6000 5024
rect 6052 4972 6058 5024
rect 6730 4972 6736 5024
rect 6788 4972 6794 5024
rect 1104 4922 8924 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 8924 4922
rect 1104 4848 8924 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 1670 4808 1676 4820
rect 1443 4780 1676 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 4617 4811 4675 4817
rect 4617 4777 4629 4811
rect 4663 4808 4675 4811
rect 4890 4808 4896 4820
rect 4663 4780 4896 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5629 4811 5687 4817
rect 5031 4780 5396 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5368 4752 5396 4780
rect 5629 4777 5641 4811
rect 5675 4808 5687 4811
rect 5994 4808 6000 4820
rect 5675 4780 6000 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6546 4768 6552 4820
rect 6604 4768 6610 4820
rect 7098 4768 7104 4820
rect 7156 4768 7162 4820
rect 8570 4768 8576 4820
rect 8628 4768 8634 4820
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 5077 4743 5135 4749
rect 5077 4740 5089 4743
rect 4764 4712 5089 4740
rect 4764 4700 4770 4712
rect 5077 4709 5089 4712
rect 5123 4709 5135 4743
rect 5077 4703 5135 4709
rect 5350 4700 5356 4752
rect 5408 4700 5414 4752
rect 6564 4740 6592 4768
rect 5736 4712 6592 4740
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 4080 4644 4353 4672
rect 2498 4564 2504 4616
rect 2556 4613 2562 4616
rect 2556 4604 2568 4613
rect 2556 4576 2601 4604
rect 2556 4567 2568 4576
rect 2556 4564 2562 4567
rect 2774 4564 2780 4616
rect 2832 4564 2838 4616
rect 4080 4536 4108 4644
rect 4341 4641 4353 4644
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 4816 4644 5672 4672
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4709 4607 4767 4613
rect 4479 4601 4660 4604
rect 4709 4601 4721 4607
rect 4479 4576 4721 4601
rect 4479 4573 4491 4576
rect 4632 4573 4721 4576
rect 4755 4604 4767 4607
rect 4816 4604 4844 4644
rect 5644 4616 5672 4644
rect 4755 4576 4844 4604
rect 4755 4573 4767 4576
rect 4433 4567 4491 4573
rect 4709 4567 4767 4573
rect 4264 4536 4292 4567
rect 4890 4564 4896 4616
rect 4948 4564 4954 4616
rect 5166 4564 5172 4616
rect 5224 4564 5230 4616
rect 5350 4564 5356 4616
rect 5408 4564 5414 4616
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 5626 4564 5632 4616
rect 5684 4564 5690 4616
rect 5736 4613 5764 4712
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 7116 4672 7144 4768
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 5960 4644 6868 4672
rect 7116 4644 7205 4672
rect 5960 4632 5966 4644
rect 6840 4616 6868 4644
rect 7193 4641 7205 4644
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6420 4576 6469 4604
rect 6420 4564 6426 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6638 4564 6644 4616
rect 6696 4564 6702 4616
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 5368 4536 5396 4564
rect 4080 4508 4200 4536
rect 4264 4508 5396 4536
rect 4172 4468 4200 4508
rect 4890 4468 4896 4480
rect 4172 4440 4896 4468
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5810 4468 5816 4480
rect 5491 4440 5816 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5810 4428 5816 4440
rect 5868 4468 5874 4480
rect 6380 4468 6408 4564
rect 6748 4536 6776 4567
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 6932 4536 6960 4564
rect 6748 4508 6960 4536
rect 7101 4539 7159 4545
rect 7101 4505 7113 4539
rect 7147 4536 7159 4539
rect 7438 4539 7496 4545
rect 7438 4536 7450 4539
rect 7147 4508 7450 4536
rect 7147 4505 7159 4508
rect 7101 4499 7159 4505
rect 7438 4505 7450 4508
rect 7484 4505 7496 4539
rect 7438 4499 7496 4505
rect 5868 4440 6408 4468
rect 5868 4428 5874 4440
rect 1104 4378 8924 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8924 4378
rect 1104 4304 8924 4326
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 4890 4264 4896 4276
rect 4764 4236 4896 4264
rect 4764 4224 4770 4236
rect 4890 4224 4896 4236
rect 4948 4264 4954 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 4948 4236 4997 4264
rect 4948 4224 4954 4236
rect 4985 4233 4997 4236
rect 5031 4233 5043 4267
rect 5442 4264 5448 4276
rect 4985 4227 5043 4233
rect 5092 4236 5448 4264
rect 4525 4199 4583 4205
rect 4525 4165 4537 4199
rect 4571 4196 4583 4199
rect 4614 4196 4620 4208
rect 4571 4168 4620 4196
rect 4571 4165 4583 4168
rect 4525 4159 4583 4165
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3234 4128 3240 4140
rect 3191 4100 3240 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 4724 4128 4752 4224
rect 3467 4100 4752 4128
rect 4985 4131 5043 4137
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 4985 4097 4997 4131
rect 5031 4097 5043 4131
rect 5092 4128 5120 4236
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 6549 4267 6607 4273
rect 6549 4233 6561 4267
rect 6595 4264 6607 4267
rect 6638 4264 6644 4276
rect 6595 4236 6644 4264
rect 6595 4233 6607 4236
rect 6549 4227 6607 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 5350 4156 5356 4208
rect 5408 4156 5414 4208
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 5092 4100 5181 4128
rect 4985 4091 5043 4097
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 3142 3884 3148 3936
rect 3200 3884 3206 3936
rect 3344 3924 3372 4091
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 5000 4060 5028 4091
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5810 4128 5816 4140
rect 5491 4100 5816 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6656 4100 6929 4128
rect 6656 4072 6684 4100
rect 6917 4097 6929 4100
rect 6963 4128 6975 4131
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 6963 4100 7205 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 7423 4100 8493 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 8481 4097 8493 4100
rect 8527 4128 8539 4131
rect 8570 4128 8576 4140
rect 8527 4100 8576 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 4212 4032 5028 4060
rect 4212 4020 4218 4032
rect 6086 4020 6092 4072
rect 6144 4020 6150 4072
rect 6638 4020 6644 4072
rect 6696 4020 6702 4072
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7055 4032 7849 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 4341 3995 4399 4001
rect 4341 3961 4353 3995
rect 4387 3992 4399 3995
rect 4706 3992 4712 4004
rect 4387 3964 4712 3992
rect 4387 3961 4399 3964
rect 4341 3955 4399 3961
rect 4706 3952 4712 3964
rect 4764 3952 4770 4004
rect 4893 3995 4951 4001
rect 4893 3961 4905 3995
rect 4939 3992 4951 3995
rect 5626 3992 5632 4004
rect 4939 3964 5632 3992
rect 4939 3961 4951 3964
rect 4893 3955 4951 3961
rect 5626 3952 5632 3964
rect 5684 3992 5690 4004
rect 6104 3992 6132 4020
rect 6840 3992 6868 4023
rect 5684 3964 6868 3992
rect 5684 3952 5690 3964
rect 3786 3924 3792 3936
rect 3344 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4522 3924 4528 3936
rect 4028 3896 4528 3924
rect 4028 3884 4034 3896
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 7285 3927 7343 3933
rect 7285 3924 7297 3927
rect 6880 3896 7297 3924
rect 6880 3884 6886 3896
rect 7285 3893 7297 3896
rect 7331 3893 7343 3927
rect 7285 3887 7343 3893
rect 1104 3834 8924 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 8924 3834
rect 1104 3760 8924 3782
rect 3142 3680 3148 3732
rect 3200 3680 3206 3732
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 3973 3723 4031 3729
rect 3973 3720 3985 3723
rect 3292 3692 3985 3720
rect 3292 3680 3298 3692
rect 3973 3689 3985 3692
rect 4019 3689 4031 3723
rect 3973 3683 4031 3689
rect 4890 3680 4896 3732
rect 4948 3680 4954 3732
rect 3160 3584 3188 3680
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4908 3652 4936 3680
rect 3927 3624 4936 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 8478 3612 8484 3664
rect 8536 3612 8542 3664
rect 3513 3587 3571 3593
rect 3513 3584 3525 3587
rect 3160 3556 3525 3584
rect 3513 3553 3525 3556
rect 3559 3553 3571 3587
rect 3513 3547 3571 3553
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 4028 3556 4077 3584
rect 4028 3544 4034 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4065 3547 4123 3553
rect 6089 3587 6147 3593
rect 6089 3553 6101 3587
rect 6135 3584 6147 3587
rect 7098 3584 7104 3596
rect 6135 3556 7104 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 3786 3476 3792 3528
rect 3844 3476 3850 3528
rect 4341 3519 4399 3525
rect 4341 3485 4353 3519
rect 4387 3516 4399 3519
rect 4798 3516 4804 3528
rect 4387 3488 4804 3516
rect 4387 3485 4399 3488
rect 4341 3479 4399 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 6638 3476 6644 3528
rect 6696 3516 6702 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 6696 3488 8309 3516
rect 6696 3476 6702 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 3804 3448 3832 3476
rect 5718 3448 5724 3460
rect 3804 3420 5724 3448
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2648 3352 2973 3380
rect 2648 3340 2654 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 1104 3290 8924 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8924 3290
rect 1104 3216 8924 3238
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4522 3176 4528 3188
rect 4387 3148 4528 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 7098 3176 7104 3188
rect 4632 3148 7104 3176
rect 2774 3108 2780 3120
rect 2332 3080 2780 3108
rect 2332 3049 2360 3080
rect 2774 3068 2780 3080
rect 2832 3108 2838 3120
rect 4632 3108 4660 3148
rect 4706 3117 4712 3120
rect 2832 3080 4660 3108
rect 2832 3068 2838 3080
rect 2590 3049 2596 3052
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2584 3040 2596 3049
rect 2551 3012 2596 3040
rect 2317 3003 2375 3009
rect 2584 3003 2596 3012
rect 2590 3000 2596 3003
rect 2648 3000 2654 3052
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4632 3040 4660 3080
rect 4700 3071 4712 3117
rect 4764 3108 4770 3120
rect 5905 3111 5963 3117
rect 4764 3080 4800 3108
rect 4706 3068 4712 3071
rect 4764 3068 4770 3080
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 5951 3080 6316 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 4479 3012 4660 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 5074 3000 5080 3052
rect 5132 3040 5138 3052
rect 6086 3040 6092 3052
rect 5132 3012 6092 3040
rect 5132 3000 5138 3012
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 6288 3040 6316 3080
rect 6362 3068 6368 3120
rect 6420 3068 6426 3120
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 6565 3111 6623 3117
rect 6565 3108 6577 3111
rect 6512 3080 6577 3108
rect 6512 3068 6518 3080
rect 6565 3077 6577 3080
rect 6611 3077 6623 3111
rect 6565 3071 6623 3077
rect 6730 3040 6736 3052
rect 6288 3012 6736 3040
rect 6181 3003 6239 3009
rect 3878 2932 3884 2984
rect 3936 2932 3942 2984
rect 3973 2975 4031 2981
rect 3973 2941 3985 2975
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 3988 2904 4016 2935
rect 4062 2932 4068 2984
rect 4120 2932 4126 2984
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2941 4215 2975
rect 6196 2972 6224 3003
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 6840 3049 6868 3148
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 7081 3043 7139 3049
rect 7081 3040 7093 3043
rect 6825 3003 6883 3009
rect 6932 3012 7093 3040
rect 6638 2972 6644 2984
rect 6196 2944 6644 2972
rect 4157 2935 4215 2941
rect 3712 2876 4016 2904
rect 3712 2848 3740 2876
rect 3694 2796 3700 2848
rect 3752 2796 3758 2848
rect 4172 2836 4200 2935
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 6932 2972 6960 3012
rect 7081 3009 7093 3012
rect 7127 3009 7139 3043
rect 7081 3003 7139 3009
rect 6748 2944 6960 2972
rect 5442 2836 5448 2848
rect 4172 2808 5448 2836
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 5810 2796 5816 2848
rect 5868 2796 5874 2848
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6227 2808 6561 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 6656 2836 6684 2932
rect 6748 2913 6776 2944
rect 6733 2907 6791 2913
rect 6733 2873 6745 2907
rect 6779 2873 6791 2907
rect 6733 2867 6791 2873
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 6656 2808 8217 2836
rect 6549 2799 6607 2805
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 1104 2746 8924 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 8924 2746
rect 1104 2672 8924 2694
rect 1489 2635 1547 2641
rect 1489 2601 1501 2635
rect 1535 2632 1547 2635
rect 1762 2632 1768 2644
rect 1535 2604 1768 2632
rect 1535 2601 1547 2604
rect 1489 2595 1547 2601
rect 1762 2592 1768 2604
rect 1820 2632 1826 2644
rect 4062 2632 4068 2644
rect 1820 2604 4068 2632
rect 1820 2592 1826 2604
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3252 2437 3280 2604
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 5074 2592 5080 2644
rect 5132 2592 5138 2644
rect 5718 2592 5724 2644
rect 5776 2592 5782 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6454 2632 6460 2644
rect 6411 2604 6460 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 4479 2468 5672 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2832 2400 2881 2428
rect 2832 2388 2838 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3510 2388 3516 2440
rect 3568 2388 3574 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 3694 2428 3700 2440
rect 3651 2400 3700 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 3694 2388 3700 2400
rect 3752 2428 3758 2440
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 3752 2400 3893 2428
rect 3752 2388 3758 2400
rect 3881 2397 3893 2400
rect 3927 2397 3939 2431
rect 3881 2391 3939 2397
rect 2624 2363 2682 2369
rect 2624 2329 2636 2363
rect 2670 2360 2682 2363
rect 3528 2360 3556 2388
rect 2670 2332 3556 2360
rect 3896 2360 3924 2391
rect 3970 2388 3976 2440
rect 4028 2428 4034 2440
rect 5644 2437 5672 2468
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 4028 2400 4537 2428
rect 4028 2388 4034 2400
rect 4525 2397 4537 2400
rect 4571 2428 4583 2431
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 4571 2400 5549 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 4709 2363 4767 2369
rect 4709 2360 4721 2363
rect 3896 2332 4721 2360
rect 2670 2329 2682 2332
rect 2624 2323 2682 2329
rect 4709 2329 4721 2332
rect 4755 2360 4767 2363
rect 5166 2360 5172 2372
rect 4755 2332 5172 2360
rect 4755 2329 4767 2332
rect 4709 2323 4767 2329
rect 5166 2320 5172 2332
rect 5224 2320 5230 2372
rect 5442 2360 5448 2372
rect 5285 2332 5448 2360
rect 2498 2252 2504 2304
rect 2556 2292 2562 2304
rect 3053 2295 3111 2301
rect 3053 2292 3065 2295
rect 2556 2264 3065 2292
rect 2556 2252 2562 2264
rect 3053 2261 3065 2264
rect 3099 2261 3111 2295
rect 3053 2255 3111 2261
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 3878 2292 3884 2304
rect 3467 2264 3884 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 4120 2264 4813 2292
rect 4120 2252 4126 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2292 4951 2295
rect 5285 2292 5313 2332
rect 5442 2320 5448 2332
rect 5500 2320 5506 2372
rect 5552 2360 5580 2391
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 6086 2388 6092 2440
rect 6144 2388 6150 2440
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6638 2428 6644 2440
rect 6595 2400 6644 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6788 2400 6837 2428
rect 6788 2388 6794 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 5828 2360 5856 2388
rect 5552 2332 5856 2360
rect 4939 2264 5313 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 5350 2252 5356 2304
rect 5408 2252 5414 2304
rect 6104 2292 6132 2388
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6104 2264 6745 2292
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 1104 2202 8924 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8924 2202
rect 1104 2128 8924 2150
<< via1 >>
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5816 9596 5868 9648
rect 6184 9528 6236 9580
rect 7288 9460 7340 9512
rect 6368 9367 6420 9376
rect 6368 9333 6377 9367
rect 6377 9333 6411 9367
rect 6411 9333 6420 9367
rect 6368 9324 6420 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2136 8916 2188 8968
rect 5724 8916 5776 8968
rect 3884 8848 3936 8900
rect 4712 8891 4764 8900
rect 4712 8857 4746 8891
rect 4746 8857 4764 8891
rect 4712 8848 4764 8857
rect 2596 8780 2648 8832
rect 5264 8780 5316 8832
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 5908 8780 5960 8832
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2136 8576 2188 8628
rect 3884 8619 3936 8628
rect 3884 8585 3893 8619
rect 3893 8585 3927 8619
rect 3927 8585 3936 8619
rect 3884 8576 3936 8585
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 5540 8508 5592 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1676 8483 1728 8492
rect 1676 8449 1710 8483
rect 1710 8449 1728 8483
rect 1676 8440 1728 8449
rect 3148 8440 3200 8492
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 5632 8440 5684 8492
rect 6920 8508 6972 8560
rect 7012 8440 7064 8492
rect 4620 8372 4672 8424
rect 2320 8236 2372 8288
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 5908 8304 5960 8356
rect 4068 8236 4120 8288
rect 4896 8236 4948 8288
rect 7288 8236 7340 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1676 8032 1728 8084
rect 2964 8032 3016 8084
rect 3240 8032 3292 8084
rect 4252 8032 4304 8084
rect 4620 8032 4672 8084
rect 4712 8032 4764 8084
rect 2596 7964 2648 8016
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 2044 7828 2096 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 3056 7828 3108 7880
rect 4528 7896 4580 7948
rect 5172 8032 5224 8084
rect 7012 8032 7064 8084
rect 3148 7760 3200 7812
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 4712 7828 4764 7880
rect 5264 7896 5316 7948
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 5724 7896 5776 7948
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 6368 7828 6420 7880
rect 7012 7828 7064 7880
rect 3976 7692 4028 7744
rect 6184 7760 6236 7812
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1768 7488 1820 7540
rect 2044 7488 2096 7540
rect 1216 7420 1268 7472
rect 2780 7420 2832 7472
rect 3056 7420 3108 7472
rect 3516 7488 3568 7540
rect 4068 7463 4120 7472
rect 4068 7429 4077 7463
rect 4077 7429 4111 7463
rect 4111 7429 4120 7463
rect 4068 7420 4120 7429
rect 4252 7420 4304 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2596 7352 2648 7404
rect 4712 7420 4764 7472
rect 5448 7488 5500 7540
rect 4528 7352 4580 7404
rect 5908 7352 5960 7404
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 1952 7284 2004 7336
rect 2688 7284 2740 7336
rect 5356 7284 5408 7336
rect 6920 7352 6972 7404
rect 6644 7284 6696 7336
rect 3700 7191 3752 7200
rect 3700 7157 3709 7191
rect 3709 7157 3743 7191
rect 3743 7157 3752 7191
rect 3700 7148 3752 7157
rect 3792 7148 3844 7200
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 7104 7352 7156 7404
rect 7196 7148 7248 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2596 6944 2648 6996
rect 3148 6987 3200 6996
rect 3148 6953 3157 6987
rect 3157 6953 3191 6987
rect 3191 6953 3200 6987
rect 3148 6944 3200 6953
rect 3792 6944 3844 6996
rect 3976 6944 4028 6996
rect 2688 6876 2740 6928
rect 1400 6808 1452 6860
rect 6460 6876 6512 6928
rect 7012 6876 7064 6928
rect 3424 6740 3476 6792
rect 1860 6715 1912 6724
rect 1860 6681 1894 6715
rect 1894 6681 1912 6715
rect 1860 6672 1912 6681
rect 5264 6715 5316 6724
rect 5264 6681 5282 6715
rect 5282 6681 5316 6715
rect 5264 6672 5316 6681
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6644 6740 6696 6792
rect 6828 6715 6880 6724
rect 6828 6681 6837 6715
rect 6837 6681 6871 6715
rect 6871 6681 6880 6715
rect 6828 6672 6880 6681
rect 5540 6604 5592 6656
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7196 6851 7248 6860
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 7288 6740 7340 6792
rect 8392 6740 8444 6792
rect 7196 6672 7248 6724
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1860 6400 1912 6452
rect 2596 6400 2648 6452
rect 3424 6400 3476 6452
rect 5264 6400 5316 6452
rect 6092 6400 6144 6452
rect 6736 6400 6788 6452
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2688 6264 2740 6316
rect 3700 6375 3752 6384
rect 3700 6341 3734 6375
rect 3734 6341 3752 6375
rect 3700 6332 3752 6341
rect 2228 6196 2280 6248
rect 4712 6264 4764 6316
rect 5080 6264 5132 6316
rect 5724 6332 5776 6384
rect 5448 6264 5500 6316
rect 5356 6128 5408 6180
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 1860 6060 1912 6112
rect 2780 6060 2832 6112
rect 3148 6060 3200 6112
rect 4712 6060 4764 6112
rect 6920 6332 6972 6384
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 6644 6196 6696 6248
rect 7104 6196 7156 6248
rect 8392 6264 8444 6316
rect 8484 6171 8536 6180
rect 8484 6137 8493 6171
rect 8493 6137 8527 6171
rect 8527 6137 8536 6171
rect 8484 6128 8536 6137
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1584 5856 1636 5908
rect 4804 5856 4856 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 7288 5856 7340 5908
rect 8576 5856 8628 5908
rect 2136 5788 2188 5840
rect 5080 5788 5132 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1860 5720 1912 5772
rect 1768 5695 1820 5704
rect 1768 5661 1778 5695
rect 1778 5661 1812 5695
rect 1812 5661 1820 5695
rect 1768 5652 1820 5661
rect 2320 5652 2372 5704
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3148 5695 3200 5704
rect 3148 5661 3157 5695
rect 3157 5661 3191 5695
rect 3191 5661 3200 5695
rect 3148 5652 3200 5661
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4620 5652 4672 5704
rect 6276 5720 6328 5772
rect 6552 5695 6604 5704
rect 6552 5661 6561 5695
rect 6561 5661 6595 5695
rect 6595 5661 6604 5695
rect 6552 5652 6604 5661
rect 2044 5627 2096 5636
rect 2044 5593 2053 5627
rect 2053 5593 2087 5627
rect 2087 5593 2096 5627
rect 2044 5584 2096 5593
rect 5356 5584 5408 5636
rect 1952 5516 2004 5568
rect 2136 5516 2188 5568
rect 2504 5516 2556 5568
rect 2596 5559 2648 5568
rect 2596 5525 2621 5559
rect 2621 5525 2648 5559
rect 2596 5516 2648 5525
rect 2780 5559 2832 5568
rect 2780 5525 2789 5559
rect 2789 5525 2823 5559
rect 2823 5525 2832 5559
rect 2780 5516 2832 5525
rect 4712 5516 4764 5568
rect 5632 5516 5684 5568
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 8576 5584 8628 5636
rect 7104 5516 7156 5568
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2044 5312 2096 5364
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 2596 5312 2648 5364
rect 2780 5244 2832 5296
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 4712 5244 4764 5296
rect 5172 5244 5224 5296
rect 5632 5287 5684 5296
rect 5632 5253 5641 5287
rect 5641 5253 5675 5287
rect 5675 5253 5684 5287
rect 5632 5244 5684 5253
rect 5816 5287 5868 5296
rect 5816 5253 5825 5287
rect 5825 5253 5859 5287
rect 5859 5253 5868 5287
rect 5816 5244 5868 5253
rect 6552 5287 6604 5296
rect 6552 5253 6561 5287
rect 6561 5253 6595 5287
rect 6595 5253 6604 5287
rect 6552 5244 6604 5253
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 7104 5312 7156 5364
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 1676 5219 1728 5228
rect 1676 5185 1685 5219
rect 1685 5185 1719 5219
rect 1719 5185 1728 5219
rect 1676 5176 1728 5185
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 5264 5176 5316 5228
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5540 5176 5592 5228
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 4988 5108 5040 5160
rect 5908 5108 5960 5160
rect 3516 5040 3568 5092
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 2780 4972 2832 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6736 4972 6788 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 1676 4768 1728 4820
rect 4896 4768 4948 4820
rect 6000 4768 6052 4820
rect 6552 4768 6604 4820
rect 7104 4768 7156 4820
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 4712 4700 4764 4752
rect 5356 4700 5408 4752
rect 2504 4607 2556 4616
rect 2504 4573 2522 4607
rect 2522 4573 2556 4607
rect 2504 4564 2556 4573
rect 2780 4607 2832 4616
rect 2780 4573 2789 4607
rect 2789 4573 2823 4607
rect 2823 4573 2832 4607
rect 2780 4564 2832 4573
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 5356 4564 5408 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 5632 4564 5684 4616
rect 5908 4632 5960 4684
rect 6368 4564 6420 4616
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 4896 4428 4948 4480
rect 5816 4428 5868 4480
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 6920 4564 6972 4616
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4712 4224 4764 4276
rect 4896 4224 4948 4276
rect 4620 4156 4672 4208
rect 3240 4088 3292 4140
rect 5448 4224 5500 4276
rect 6644 4224 6696 4276
rect 5356 4199 5408 4208
rect 5356 4165 5365 4199
rect 5365 4165 5399 4199
rect 5399 4165 5408 4199
rect 5356 4156 5408 4165
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 4160 4020 4212 4072
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5816 4088 5868 4140
rect 8576 4088 8628 4140
rect 6092 4020 6144 4072
rect 6644 4020 6696 4072
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 4712 3952 4764 4004
rect 5632 3952 5684 4004
rect 3792 3884 3844 3936
rect 3976 3884 4028 3936
rect 4528 3927 4580 3936
rect 4528 3893 4537 3927
rect 4537 3893 4571 3927
rect 4571 3893 4580 3927
rect 4528 3884 4580 3893
rect 6828 3884 6880 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3148 3680 3200 3732
rect 3240 3680 3292 3732
rect 4896 3680 4948 3732
rect 8484 3655 8536 3664
rect 8484 3621 8493 3655
rect 8493 3621 8527 3655
rect 8527 3621 8536 3655
rect 8484 3612 8536 3621
rect 3976 3544 4028 3596
rect 7104 3544 7156 3596
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 4804 3476 4856 3528
rect 6644 3476 6696 3528
rect 5724 3408 5776 3460
rect 2596 3340 2648 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4528 3136 4580 3188
rect 2780 3068 2832 3120
rect 2596 3043 2648 3052
rect 2596 3009 2630 3043
rect 2630 3009 2648 3043
rect 2596 3000 2648 3009
rect 4712 3111 4764 3120
rect 4712 3077 4746 3111
rect 4746 3077 4764 3111
rect 4712 3068 4764 3077
rect 5080 3000 5132 3052
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 6368 3111 6420 3120
rect 6368 3077 6377 3111
rect 6377 3077 6411 3111
rect 6411 3077 6420 3111
rect 6368 3068 6420 3077
rect 6460 3068 6512 3120
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 6736 3000 6788 3052
rect 7104 3136 7156 3188
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 6644 2932 6696 2984
rect 5448 2796 5500 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 1768 2592 1820 2644
rect 2780 2388 2832 2440
rect 4068 2592 4120 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 6460 2592 6512 2644
rect 3516 2388 3568 2440
rect 3700 2388 3752 2440
rect 3976 2388 4028 2440
rect 5172 2320 5224 2372
rect 2504 2252 2556 2304
rect 3884 2252 3936 2304
rect 4068 2252 4120 2304
rect 5448 2320 5500 2372
rect 5816 2388 5868 2440
rect 6092 2388 6144 2440
rect 6644 2388 6696 2440
rect 6736 2388 6788 2440
rect 5356 2295 5408 2304
rect 5356 2261 5365 2295
rect 5365 2261 5399 2295
rect 5399 2261 5408 2295
rect 5356 2252 5408 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5814 11398 5870 12198
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5828 9654 5856 11398
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 2148 8634 2176 8910
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1214 7576 1270 7585
rect 1214 7511 1270 7520
rect 1228 7478 1256 7511
rect 1216 7472 1268 7478
rect 1216 7414 1268 7420
rect 1412 6866 1440 8434
rect 1688 8090 1716 8434
rect 2320 8288 2372 8294
rect 2240 8248 2320 8276
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 1780 7546 1808 7822
rect 2056 7546 2084 7822
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6458 1900 6666
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1676 6316 1728 6322
rect 1412 5710 1440 6287
rect 1676 6258 1728 6264
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1504 4865 1532 6054
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1596 5234 1624 5850
rect 1688 5234 1716 6258
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5778 1900 6054
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1490 4856 1546 4865
rect 1688 4826 1716 5170
rect 1490 4791 1546 4800
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1780 2650 1808 5646
rect 1964 5574 1992 7278
rect 2056 6322 2084 7482
rect 2240 7410 2268 8248
rect 2320 8230 2372 8236
rect 2608 8022 2636 8774
rect 3896 8634 3924 8842
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3160 8378 3188 8434
rect 3068 8350 3188 8378
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 8090 3004 8230
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2596 8016 2648 8022
rect 2648 7964 2728 7970
rect 2596 7958 2728 7964
rect 2608 7942 2728 7958
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2608 7410 2636 7822
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2044 6316 2096 6322
rect 2096 6276 2176 6304
rect 2044 6258 2096 6264
rect 2148 5846 2176 6276
rect 2240 6254 2268 7346
rect 2608 7002 2636 7346
rect 2700 7342 2728 7942
rect 3068 7886 3096 8350
rect 3252 8090 3280 8434
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7478 3096 7822
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2608 6458 2636 6938
rect 2700 6934 2728 7278
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2700 6322 2728 6870
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2792 6118 2820 7414
rect 3160 7002 3188 7754
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3528 7546 3556 7686
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3436 6458 3464 6734
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3712 6390 3740 7142
rect 3804 7002 3832 7142
rect 3988 7002 4016 7686
rect 4080 7478 4108 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 8366
rect 4724 8090 4752 8842
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4264 7478 4292 8026
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4068 7472 4120 7478
rect 4068 7414 4120 7420
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4540 7410 4568 7890
rect 4712 7880 4764 7886
rect 4618 7848 4674 7857
rect 4908 7868 4936 8230
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5184 7886 5212 8026
rect 5276 7954 5304 8774
rect 5736 8634 5764 8910
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5552 7886 5580 8502
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 4764 7840 4936 7868
rect 5172 7880 5224 7886
rect 4712 7822 4764 7828
rect 5172 7822 5224 7828
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 4618 7783 4674 7792
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3700 6384 3752 6390
rect 3700 6326 3752 6332
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 2044 5636 2096 5642
rect 2044 5578 2096 5584
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 2056 5370 2084 5578
rect 2148 5574 2176 5782
rect 3160 5710 3188 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5710 4660 7783
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5460 7546 5488 7822
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4724 6322 4752 7414
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5264 6724 5316 6730
rect 5264 6666 5316 6672
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6458 5304 6666
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 2332 5370 2360 5646
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2780 5568 2832 5574
rect 3068 5545 3096 5646
rect 2780 5510 2832 5516
rect 3054 5536 3110 5545
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2516 4622 2544 5510
rect 2608 5370 2636 5510
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2792 5302 2820 5510
rect 3054 5471 3110 5480
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 4080 5234 4108 5646
rect 4724 5574 4752 6054
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 5302 4752 5510
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4622 2820 4966
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2608 3058 2636 3334
rect 2792 3126 2820 4558
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 3738 3188 3878
rect 3252 3738 3280 4082
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 2792 2446 2820 3062
rect 3528 2446 3556 5034
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4724 4842 4752 5238
rect 4632 4814 4752 4842
rect 4632 4706 4660 4814
rect 4540 4678 4660 4706
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4172 4078 4200 4558
rect 4160 4072 4212 4078
rect 4080 4020 4160 4026
rect 4080 4014 4212 4020
rect 4080 3998 4200 4014
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3804 3534 3832 3878
rect 3988 3602 4016 3878
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 4080 2990 4108 3998
rect 4540 3942 4568 4678
rect 4724 4282 4752 4694
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3210 4660 4150
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4540 3194 4660 3210
rect 4528 3188 4660 3194
rect 4580 3182 4660 3188
rect 4528 3130 4580 3136
rect 4724 3126 4752 3946
rect 4816 3534 4844 5850
rect 5092 5846 5120 6258
rect 5368 6186 5396 7278
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6322 5488 7142
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5356 6180 5408 6186
rect 5408 6140 5488 6168
rect 5356 6122 5408 6128
rect 5080 5840 5132 5846
rect 5132 5800 5304 5828
rect 5080 5782 5132 5788
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4826 4936 4966
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5000 4706 5028 5102
rect 4908 4678 5028 4706
rect 4908 4622 4936 4678
rect 5184 4622 5212 5238
rect 5276 5234 5304 5800
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5370 5396 5578
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5368 4758 5396 5170
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5368 4622 5396 4694
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4908 4486 4936 4558
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4908 3738 4936 4218
rect 5368 4214 5396 4558
rect 5460 4282 5488 6140
rect 5552 5234 5580 6598
rect 5644 5914 5672 8434
rect 5920 8362 5948 8774
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5736 6390 5764 7890
rect 5920 7410 5948 8298
rect 6196 7818 6224 9522
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 7886 6408 9318
rect 7300 8974 7328 9454
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6184 7812 6236 7818
rect 6184 7754 6236 7760
rect 6196 7410 6224 7754
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6656 7342 6684 8774
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6932 7410 6960 8502
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7024 8090 7052 8434
rect 7300 8294 7328 8910
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 7024 6934 7052 7822
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 6472 6798 6500 6870
rect 7024 6798 7052 6870
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6104 6458 6132 6598
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 6288 5778 6316 6734
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6472 5692 6500 6734
rect 6656 6254 6684 6734
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6458 6776 6598
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6552 5704 6604 5710
rect 6472 5664 6552 5692
rect 6552 5646 6604 5652
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5644 5302 5672 5510
rect 6564 5302 6592 5646
rect 6644 5568 6696 5574
rect 6696 5528 6776 5556
rect 6644 5510 6696 5516
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5552 4622 5580 5170
rect 5644 4622 5672 5238
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5552 4468 5580 4558
rect 5828 4486 5856 5238
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4690 5948 5102
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4826 6040 4966
rect 6564 4826 6592 5238
rect 6748 5030 6776 5528
rect 6840 5234 6868 6666
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6932 5370 6960 6326
rect 7116 6254 7144 7346
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 7208 6866 7236 7142
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 8404 6798 8432 7142
rect 8496 6905 8524 7686
rect 8482 6896 8538 6905
rect 8482 6831 8538 6840
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7208 6458 7236 6666
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7300 5914 7328 6734
rect 8404 6322 8432 6734
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8482 6216 8538 6225
rect 8482 6151 8484 6160
rect 8536 6151 8538 6160
rect 8484 6122 8536 6128
rect 8588 5914 8616 6598
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 8116 5568 8168 5574
rect 8484 5568 8536 5574
rect 8116 5510 8168 5516
rect 8482 5536 8484 5545
rect 8536 5536 8538 5545
rect 7116 5370 7144 5510
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 5816 4480 5868 4486
rect 5552 4440 5672 4468
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2446 3740 2790
rect 3896 2774 3924 2926
rect 3896 2746 4016 2774
rect 3988 2446 4016 2746
rect 4080 2650 4108 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5092 2650 5120 2994
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4080 2310 4108 2586
rect 5172 2372 5224 2378
rect 5276 2360 5304 4082
rect 5460 2854 5488 4218
rect 5644 4010 5672 4440
rect 5816 4422 5868 4428
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2378 5488 2790
rect 5736 2650 5764 3402
rect 5828 2854 5856 4082
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6104 3058 6132 4014
rect 6380 3126 6408 4558
rect 6656 4282 6684 4558
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6748 4078 6776 4966
rect 6932 4622 6960 5306
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 4826 7144 5102
rect 8128 4865 8156 5510
rect 8482 5471 8538 5480
rect 8114 4856 8170 4865
rect 7104 4820 7156 4826
rect 8588 4826 8616 5578
rect 8114 4791 8170 4800
rect 8576 4820 8628 4826
rect 7104 4762 7156 4768
rect 8576 4762 8628 4768
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6656 3534 6684 4014
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5828 2446 5856 2790
rect 6104 2446 6132 2994
rect 6472 2650 6500 3062
rect 6656 2990 6684 3470
rect 6748 3058 6776 4014
rect 6840 3942 6868 4558
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 7116 3602 7144 4762
rect 8588 4146 8616 4762
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 3194 7144 3538
rect 8496 3505 8524 3606
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6656 2446 6684 2926
rect 6748 2446 6776 2994
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 5224 2332 5304 2360
rect 5448 2372 5500 2378
rect 5172 2314 5224 2320
rect 5448 2314 5500 2320
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 2516 1170 2544 2246
rect 2516 1142 2636 1170
rect 2608 800 2636 1142
rect 3896 800 3924 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5368 1170 5396 2246
rect 5184 1142 5396 1170
rect 5184 800 5212 1142
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
<< via2 >>
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1214 7520 1270 7576
rect 1398 6296 1454 6352
rect 1490 4800 1546 4856
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4618 7792 4674 7848
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 3054 5480 3110 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 8482 6840 8538 6896
rect 8482 6180 8538 6216
rect 8482 6160 8484 6180
rect 8484 6160 8536 6180
rect 8536 6160 8538 6180
rect 8482 5516 8484 5536
rect 8484 5516 8536 5536
rect 8536 5516 8538 5536
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8482 5480 8538 5516
rect 8114 4800 8170 4856
rect 8482 3440 8538 3496
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 0 8198 2790 8258
rect 0 8168 800 8198
rect 2730 7850 2790 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4613 7850 4679 7853
rect 2730 7848 4679 7850
rect 2730 7792 4618 7848
rect 4674 7792 4679 7848
rect 2730 7790 4679 7792
rect 4613 7787 4679 7790
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1209 7578 1275 7581
rect 0 7488 858 7578
rect 798 7442 858 7488
rect 1166 7576 1275 7578
rect 1166 7520 1214 7576
rect 1270 7520 1275 7576
rect 1166 7515 1275 7520
rect 1166 7442 1226 7515
rect 798 7382 1226 7442
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6900 800 6928
rect 0 6836 796 6900
rect 860 6836 866 6900
rect 8477 6898 8543 6901
rect 9254 6898 10054 6928
rect 8477 6896 10054 6898
rect 8477 6840 8482 6896
rect 8538 6840 10054 6896
rect 8477 6838 10054 6840
rect 0 6808 800 6836
rect 8477 6835 8543 6838
rect 9254 6808 10054 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 790 6292 796 6356
rect 860 6354 866 6356
rect 1393 6354 1459 6357
rect 860 6352 1459 6354
rect 860 6296 1398 6352
rect 1454 6296 1459 6352
rect 860 6294 1459 6296
rect 860 6292 866 6294
rect 1393 6291 1459 6294
rect 8477 6218 8543 6221
rect 9254 6218 10054 6248
rect 8477 6216 10054 6218
rect 8477 6160 8482 6216
rect 8538 6160 10054 6216
rect 8477 6158 10054 6160
rect 8477 6155 8543 6158
rect 9254 6128 10054 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 3049 5538 3115 5541
rect 0 5536 3115 5538
rect 0 5480 3054 5536
rect 3110 5480 3115 5536
rect 0 5478 3115 5480
rect 0 5448 800 5478
rect 3049 5475 3115 5478
rect 8477 5538 8543 5541
rect 9254 5538 10054 5568
rect 8477 5536 10054 5538
rect 8477 5480 8482 5536
rect 8538 5480 10054 5536
rect 8477 5478 10054 5480
rect 8477 5475 8543 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 9254 5448 10054 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 8109 4858 8175 4861
rect 9254 4858 10054 4888
rect 8109 4856 10054 4858
rect 8109 4800 8114 4856
rect 8170 4800 10054 4856
rect 8109 4798 10054 4800
rect 8109 4795 8175 4798
rect 9254 4768 10054 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 8477 3498 8543 3501
rect 9254 3498 10054 3528
rect 8477 3496 10054 3498
rect 8477 3440 8482 3496
rect 8538 3440 10054 3496
rect 8477 3438 10054 3440
rect 8477 3435 8543 3438
rect 9254 3408 10054 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 796 6836 860 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 796 6292 860 6356
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9840
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 795 6900 861 6901
rect 795 6836 796 6900
rect 860 6836 861 6900
rect 795 6835 861 6836
rect 798 6357 858 6835
rect 795 6356 861 6357
rect 795 6292 796 6356
rect 860 6292 861 6356
rect 795 6291 861 6292
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 9824 5188 9840
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _049_
timestamp -3599
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp -3599
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _051_
timestamp -3599
transform -1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _052_
timestamp -3599
transform 1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _053_
timestamp -3599
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _054_
timestamp -3599
transform -1 0 6624 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _055_
timestamp -3599
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _056_
timestamp -3599
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _057_
timestamp -3599
transform 1 0 5336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _058_
timestamp -3599
transform -1 0 4692 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _059_
timestamp -3599
transform -1 0 5336 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _060_
timestamp -3599
transform 1 0 1656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _061_
timestamp -3599
transform 1 0 3864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _062_
timestamp -3599
transform -1 0 5428 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _063_
timestamp -3599
transform -1 0 3128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _064_
timestamp -3599
transform -1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _065_
timestamp -3599
transform 1 0 2392 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _066_
timestamp -3599
transform -1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp -3599
transform 1 0 1840 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _068_
timestamp -3599
transform -1 0 2024 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _069_
timestamp -3599
transform 1 0 2300 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _070_
timestamp -3599
transform -1 0 2208 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _071_
timestamp -3599
transform -1 0 3680 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _072_
timestamp -3599
transform 1 0 4416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _073_
timestamp -3599
transform -1 0 5888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _074_
timestamp -3599
transform -1 0 3680 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _075_
timestamp -3599
transform -1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _076_
timestamp -3599
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _077_
timestamp -3599
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _078_
timestamp -3599
transform 1 0 3128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _079_
timestamp -3599
transform -1 0 4416 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _080_
timestamp -3599
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _081_
timestamp -3599
transform -1 0 4968 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _082_
timestamp -3599
transform -1 0 5520 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _083_
timestamp -3599
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _084_
timestamp -3599
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _085_
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _086_
timestamp -3599
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _087_
timestamp -3599
transform -1 0 6164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _088_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _089_
timestamp -3599
transform -1 0 6808 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _090_
timestamp -3599
transform -1 0 7084 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _091_
timestamp -3599
transform -1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _092_
timestamp -3599
transform 1 0 6808 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _093_
timestamp -3599
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _094_
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _095_
timestamp -3599
transform 1 0 6348 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _096_
timestamp -3599
transform 1 0 6532 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _097_
timestamp -3599
transform -1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _098_
timestamp -3599
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _099_
timestamp -3599
transform -1 0 2944 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _100_
timestamp -3599
transform 1 0 2392 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _101_
timestamp -3599
transform -1 0 3588 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _102_
timestamp -3599
transform -1 0 5612 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _103_
timestamp -3599
transform 1 0 3404 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _104_
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _105_
timestamp -3599
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _106_
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _107_
timestamp -3599
transform 1 0 4416 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp -3599
transform 1 0 2300 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _109_
timestamp -3599
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _110_
timestamp -3599
transform 1 0 7084 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _111_
timestamp -3599
transform 1 0 6992 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _112_
timestamp -3599
transform 1 0 7176 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _113_
timestamp -3599
transform 1 0 6808 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _114_
timestamp -3599
transform 1 0 7176 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 4324 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -3599
transform 1 0 4324 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -3599
transform 1 0 4416 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_52
timestamp -3599
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_63
timestamp 1636964856
transform 1 0 6900 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_75
timestamp -3599
transform 1 0 8004 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_11
timestamp -3599
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_78
timestamp -3599
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_15
timestamp -3599
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_19
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_33
timestamp -3599
transform 1 0 4140 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_55
timestamp 1636964856
transform 1 0 6164 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_67
timestamp -3599
transform 1 0 7268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_75
timestamp -3599
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp -3599
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp -3599
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_26
timestamp -3599
transform 1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_34
timestamp -3599
transform 1 0 4232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_48
timestamp -3599
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp -3599
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_69
timestamp -3599
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_81
timestamp -3599
transform 1 0 8556 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp -3599
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_29
timestamp -3599
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_51
timestamp -3599
transform 1 0 5796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_57
timestamp -3599
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_30
timestamp -3599
transform 1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_50
timestamp -3599
transform 1 0 5704 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_81
timestamp -3599
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp -3599
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_33
timestamp -3599
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_65
timestamp -3599
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_73
timestamp -3599
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_12
timestamp -3599
transform 1 0 2208 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_22
timestamp -3599
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_47
timestamp -3599
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp -3599
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_67
timestamp -3599
transform 1 0 7268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_75
timestamp -3599
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_21
timestamp -3599
transform 1 0 3036 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_7
timestamp -3599
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_17
timestamp -3599
transform 1 0 2668 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_60
timestamp -3599
transform 1 0 6624 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_80
timestamp -3599
transform 1 0 8464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_10
timestamp -3599
transform 1 0 2024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_52
timestamp -3599
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_64
timestamp 1636964856
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_76
timestamp -3599
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_22
timestamp -3599
transform 1 0 3128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_31
timestamp -3599
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_35
timestamp -3599
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_73
timestamp -3599
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_81
timestamp -3599
transform 1 0 8556 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp -3599
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp -3599
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_35
timestamp -3599
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_68
timestamp 1636964856
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_80
timestamp -3599
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636964856
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636964856
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp -3599
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 1636964856
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1636964856
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp -3599
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_71
timestamp -3599
transform 1 0 7636 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_79
timestamp -3599
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -3599
transform 1 0 4048 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -3599
transform 1 0 1656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -3599
transform 1 0 5888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -3599
transform 1 0 4784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp -3599
transform -1 0 3680 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp -3599
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp -3599
transform -1 0 6256 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp -3599
transform 1 0 6256 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp -3599
transform -1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp -3599
transform 1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp -3599
transform -1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp -3599
transform -1 0 5152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -3599
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp -3599
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform -1 0 3128 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output4
timestamp -3599
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp -3599
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp -3599
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp -3599
transform 1 0 8280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp -3599
transform 1 0 8280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -3599
transform 1 0 7912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp -3599
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp -3599
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp -3599
transform 1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 8924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 8924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 8924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_32
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_33
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_34
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_35
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_36
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_37
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_38
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_39
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_40
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_41
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_42
timestamp -3599
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_43
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 count_out[0]
port 3 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 count_out[1]
port 4 nsew signal output
flabel metal3 s 9254 6808 10054 6928 0 FreeSans 480 0 0 0 count_out[2]
port 5 nsew signal output
flabel metal3 s 9254 6128 10054 6248 0 FreeSans 480 0 0 0 count_out[3]
port 6 nsew signal output
flabel metal3 s 9254 5448 10054 5568 0 FreeSans 480 0 0 0 count_out[4]
port 7 nsew signal output
flabel metal3 s 9254 3408 10054 3528 0 FreeSans 480 0 0 0 count_out[5]
port 8 nsew signal output
flabel metal3 s 9254 4768 10054 4888 0 FreeSans 480 0 0 0 count_out[6]
port 9 nsew signal output
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 data_in
port 10 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 ready
port 11 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 rst
port 12 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 running
port 13 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 start
port 14 nsew signal input
flabel metal2 s 5814 11398 5870 12198 0 FreeSans 224 90 0 0 temp_reset
port 15 nsew signal output
rlabel via1 5014 9792 5014 9792 0 VGND
rlabel metal1 5014 9248 5014 9248 0 VPWR
rlabel metal2 2806 5406 2806 5406 0 _000_
rlabel via1 3721 6358 3721 6358 0 _001_
rlabel via1 2534 4590 2534 4590 0 _002_
rlabel metal1 3097 2346 3097 2346 0 _003_
rlabel metal2 3910 8738 3910 8738 0 _004_
rlabel metal1 5336 6426 5336 6426 0 _005_
rlabel metal1 1656 8058 1656 8058 0 _006_
rlabel metal1 1840 6426 1840 6426 0 _007_
rlabel metal1 6072 7922 6072 7922 0 _008_
rlabel metal1 3956 7990 3956 7990 0 _009_
rlabel metal1 3358 3570 3358 3570 0 _010_
rlabel via1 4733 3094 4733 3094 0 _011_
rlabel metal1 7068 5270 7068 5270 0 _012_
rlabel metal1 6854 6086 6854 6086 0 _013_
rlabel metal2 7222 6562 7222 6562 0 _014_
rlabel metal1 7028 3026 7028 3026 0 _015_
rlabel metal1 7298 4522 7298 4522 0 _016_
rlabel metal1 3818 3468 3818 3468 0 _017_
rlabel metal1 6072 7514 6072 7514 0 _018_
rlabel metal2 2990 8160 2990 8160 0 _019_
rlabel metal2 2070 7072 2070 7072 0 _020_
rlabel metal1 1794 5338 1794 5338 0 _021_
rlabel metal2 5658 5406 5658 5406 0 _022_
rlabel metal2 6854 4250 6854 4250 0 _023_
rlabel metal1 5198 4794 5198 4794 0 _024_
rlabel metal1 1978 5712 1978 5712 0 _025_
rlabel metal1 4784 4794 4784 4794 0 _026_
rlabel metal1 4462 7412 4462 7412 0 _027_
rlabel metal1 3174 8058 3174 8058 0 _028_
rlabel metal1 1840 7514 1840 7514 0 _029_
rlabel metal1 1978 6222 1978 6222 0 _030_
rlabel metal2 3174 7378 3174 7378 0 _031_
rlabel metal1 4600 7242 4600 7242 0 _032_
rlabel metal1 4876 4250 4876 4250 0 _033_
rlabel metal1 6624 6358 6624 6358 0 _034_
rlabel metal1 3634 3706 3634 3706 0 _035_
rlabel metal1 4462 3162 4462 3162 0 _036_
rlabel metal1 5612 3026 5612 3026 0 _037_
rlabel metal1 6440 4590 6440 4590 0 _038_
rlabel metal1 5842 4794 5842 4794 0 _039_
rlabel metal1 6226 5270 6226 5270 0 _040_
rlabel metal1 6624 6086 6624 6086 0 _041_
rlabel metal1 6356 6426 6356 6426 0 _042_
rlabel metal1 7130 6086 7130 6086 0 _043_
rlabel metal1 6808 2414 6808 2414 0 _044_
rlabel metal2 6946 5848 6946 5848 0 _045_
rlabel metal1 6394 2822 6394 2822 0 _046_
rlabel metal1 6440 2618 6440 2618 0 _047_
rlabel metal1 6624 4250 6624 4250 0 _048_
rlabel metal3 1717 8228 1717 8228 0 clk
rlabel metal2 5658 7174 5658 7174 0 clknet_0_clk
rlabel metal1 2852 2414 2852 2414 0 clknet_1_0__leaf_clk
rlabel metal1 1426 8500 1426 8500 0 clknet_1_1__leaf_clk
rlabel metal2 4094 5440 4094 5440 0 controller_inst.clear
rlabel metal2 3910 1520 3910 1520 0 count_out[0]
rlabel metal2 5198 959 5198 959 0 count_out[1]
rlabel metal2 8510 7293 8510 7293 0 count_out[2]
rlabel via2 8510 6171 8510 6171 0 count_out[3]
rlabel via2 8510 5525 8510 5525 0 count_out[4]
rlabel metal2 8510 3553 8510 3553 0 count_out[5]
rlabel metal2 8142 5185 8142 5185 0 count_out[6]
rlabel metal1 5106 6154 5106 6154 0 data_counter_inst.inc
rlabel metal2 2254 6800 2254 6800 0 data_edge_detector_inst.input_buffer\[0\]
rlabel metal2 2622 7616 2622 7616 0 data_edge_detector_inst.input_buffer\[1\]
rlabel metal1 6348 8262 6348 8262 0 data_edge_detector_inst.reset_counter\[0\]
rlabel metal1 5566 8806 5566 8806 0 data_edge_detector_inst.reset_counter\[1\]
rlabel metal2 2622 8398 2622 8398 0 data_edge_detector_inst.state\[0\]
rlabel metal3 751 6868 751 6868 0 data_in
rlabel metal1 1794 5542 1794 5542 0 net1
rlabel metal2 8602 5202 8602 5202 0 net10
rlabel metal2 1702 5746 1702 5746 0 net11
rlabel metal1 1656 2618 1656 2618 0 net12
rlabel metal2 6210 8466 6210 8466 0 net13
rlabel metal1 4784 5134 4784 5134 0 net14
rlabel metal1 2484 5338 2484 5338 0 net15
rlabel metal1 6256 8806 6256 8806 0 net16
rlabel metal1 5198 6222 5198 6222 0 net17
rlabel metal1 5658 2448 5658 2448 0 net18
rlabel via1 2617 3026 2617 3026 0 net19
rlabel metal2 1886 5916 1886 5916 0 net2
rlabel metal1 5980 7854 5980 7854 0 net20
rlabel metal1 5520 7514 5520 7514 0 net21
rlabel metal1 6992 8058 6992 8058 0 net22
rlabel metal1 7452 4046 7452 4046 0 net23
rlabel metal1 4002 7378 4002 7378 0 net24
rlabel metal1 4738 7276 4738 7276 0 net25
rlabel metal1 4554 8058 4554 8058 0 net26
rlabel metal1 2116 5882 2116 5882 0 net3
rlabel metal1 4968 2346 4968 2346 0 net4
rlabel metal1 5566 2380 5566 2380 0 net5
rlabel metal2 7038 7310 7038 7310 0 net6
rlabel metal1 8372 6290 8372 6290 0 net7
rlabel metal1 8464 5678 8464 5678 0 net8
rlabel metal1 6624 2414 6624 2414 0 net9
rlabel metal3 1096 4828 1096 4828 0 ready
rlabel metal3 751 7548 751 7548 0 rst
rlabel metal2 2622 959 2622 959 0 running
rlabel metal2 3082 5593 3082 5593 0 start
rlabel metal1 6716 9622 6716 9622 0 temp_reset
<< properties >>
string FIXED_BBOX 0 0 10054 12198
<< end >>

.subckt top_verilog clk rst data_in start ready running temp_reset d7 d6 d5 d4 d3 d2 d1 d0

adut [clk rst data_in start] [ready running temp_reset d7 d6 d5 d4 d3 d2 d1 d0] null top 
.model top d_cosim simulation="../../../design/time-to-digital/build/top.so" 
.ends
*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR04_lpe.spi
#else
.include ../../../work/xsch/CNR_GR04.spice
.include ../../../work/xsch/CNR_GR04_T2I_PK.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
*.param TRF = 10p

*.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc 1.8
VOUT I_OUT r01 dc 0 
R0  r01 VSS 1k

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
*.include ../xdut.spi
XDUT VDD_1V8 VSS I_OUT CNR_GR04

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------
.save all i(VDD) i(VOUT)

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save ${VPORTS}
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*optran 0 0 0 100p 2n 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
*tran 10p 10n 1p

dc TEMP -40 125 5

write
quit
#endif

.endc

.end

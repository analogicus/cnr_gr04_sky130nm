magic
tech sky130B
magscale 1 2
timestamp 1713180773
<< error_s >>
rect 3404 9096 3612 9102
rect 3404 9084 3416 9096
rect 3600 9084 3612 9096
rect 3398 7906 3414 8110
rect 3398 7884 3618 7906
rect 3630 7884 3646 8110
rect 7360 7898 7372 7904
rect 7412 7898 7424 7904
rect 7348 7880 7354 7892
rect 7430 7880 7436 7892
rect 6487 6912 6505 6918
rect 6567 6912 6585 6918
rect 6481 6894 6487 6912
rect 6585 6894 6591 6912
rect 6481 6814 6487 6832
rect 6585 6814 6591 6832
rect 6487 6808 6505 6814
rect 6567 6808 6585 6814
rect 5676 6592 5688 6598
rect 5664 6574 5670 6586
rect 5664 6522 5670 6534
rect 5686 6532 5730 6556
rect 7786 6540 7830 6556
rect 5676 6510 5688 6516
rect 5260 6304 5272 6310
rect 5248 6286 5254 6298
rect 5248 6234 5254 6246
rect 5260 6222 5272 6228
rect 6708 5652 6714 5658
rect 6766 5652 6772 5658
rect 6702 5646 6708 5652
rect 6772 5646 6778 5652
rect 6702 5588 6708 5594
rect 6772 5588 6778 5594
rect 6708 5582 6714 5588
rect 6766 5582 6772 5588
rect 5644 4904 5656 4910
rect 5632 4886 5638 4898
rect 5632 4834 5638 4846
rect 5644 4822 5656 4828
rect 4504 2091 5464 2411
rect 4765 2090 5464 2091
rect 4094 1987 4167 2015
rect 4529 1981 4547 1987
rect 4572 1981 4590 1987
rect 4523 1963 4529 1981
rect 4590 1963 4596 1981
rect 4094 1908 4167 1936
rect 4523 1920 4529 1938
rect 4590 1920 4596 1938
rect 4529 1914 4547 1920
rect 4572 1914 4590 1920
rect 4780 1771 5464 2090
rect 5728 1856 5734 2044
rect 5897 1917 5916 2044
rect 6708 2012 6726 2018
rect 6754 2012 6772 2018
rect 5935 1955 5954 2006
rect 5980 1955 5986 2006
rect 6702 1994 6708 2012
rect 6772 1994 6778 2012
rect 8324 1968 8476 2004
rect 6702 1948 6708 1966
rect 6772 1948 6778 1966
rect 8324 1956 8360 1968
rect 8440 1956 8476 1968
rect 6708 1942 6726 1948
rect 6754 1942 6772 1948
rect 8324 1940 8476 1956
rect 8324 1880 8360 1940
rect 8374 1936 8426 1940
rect 8440 1880 8476 1940
rect 8324 1844 8476 1880
rect 4780 1727 5188 1771
rect 3462 1170 3478 1176
rect 3490 1132 3506 1170
rect 3490 1110 3550 1132
<< nsubdiff >>
rect 4816 2091 5152 2099
rect 4816 1771 4824 2091
rect 5144 1771 5152 2091
rect 8360 1956 8440 1968
rect 8360 1892 8368 1956
rect 8432 1892 8440 1956
rect 8360 1880 8440 1892
rect 4816 1763 5152 1771
<< nsubdiffcont >>
rect 8368 1892 8432 1956
<< poly >>
rect 5676 6576 5740 6592
rect 5676 6532 5686 6576
rect 5730 6532 5740 6576
rect 5676 6516 5740 6532
rect 7776 6584 7840 6600
rect 7776 6540 7786 6584
rect 7830 6540 7840 6584
rect 7776 6524 7840 6540
<< polycont >>
rect 5686 6532 5730 6576
rect 7786 6540 7830 6584
<< locali >>
rect 3400 9100 3404 9300
rect 3612 9100 8200 9300
rect 6337 8628 6423 9100
rect 4637 8542 8163 8628
rect 4580 6820 6493 6906
rect 6579 6820 8236 6906
rect 4637 6666 4723 6820
rect 5977 6666 6063 6820
rect 6737 6666 6823 6820
rect 8097 6666 8183 6820
rect 5670 6532 5676 6576
rect 5740 6532 5746 6576
rect 7770 6540 7776 6584
rect 7840 6540 7846 6584
rect 7057 5357 8863 5443
rect 5740 5180 5770 5280
rect 5870 5180 5880 5280
rect 7057 5278 7143 5357
rect 8777 5297 8863 5357
rect 4630 4320 4690 4470
rect 6370 4320 6430 4470
rect 4580 4280 6500 4320
rect 5764 4260 6500 4280
rect 5728 2044 5986 2074
rect 5916 2006 5986 2044
rect 8374 2026 8426 2074
rect 5916 1955 5935 2006
rect 5916 1954 5986 1955
rect 8352 1892 8368 1956
rect 8432 1892 8448 1956
rect 3040 1825 3118 1826
rect 5728 1788 5916 1856
rect 3040 1746 3118 1747
<< viali >>
rect 3404 9096 3612 9304
rect -566 8312 -346 8532
rect 5676 8368 5740 8432
rect 7794 8374 7846 8426
rect 5260 7828 5324 7892
rect 5674 7834 5726 7886
rect 7360 7828 7424 7892
rect 6493 6820 6579 6906
rect 5334 6594 5386 6646
rect 7366 6594 7418 6646
rect 5676 6576 5740 6586
rect 7776 6584 7840 6594
rect 5676 6532 5686 6576
rect 5686 6532 5730 6576
rect 5730 6532 5740 6576
rect 7776 6540 7786 6584
rect 7786 6540 7830 6584
rect 7830 6540 7840 6584
rect 5676 6522 5740 6532
rect 7776 6530 7840 6540
rect 5260 6234 5324 6298
rect 7354 6240 7406 6292
rect 5770 5180 5870 5280
rect 6036 5116 6124 5204
rect 7374 5194 7426 5246
rect 5644 4834 5708 4898
rect 6334 4840 6386 4892
rect 6060 4548 6124 4612
rect 8454 4554 8506 4606
rect 4972 4474 5044 4546
rect 8044 4270 8108 4334
rect 8754 4276 8806 4328
rect 4535 1926 4584 1975
rect 5728 1856 5916 2044
rect 5935 1955 5986 2006
rect 6714 1954 6766 2006
rect 8374 1974 8426 2026
rect 8374 1898 8426 1950
rect 3040 1747 3118 1825
rect -442 1182 -382 1242
<< metal1 >>
rect -566 9736 3662 9956
rect -566 8538 -346 9736
rect 3442 9316 3662 9736
rect 3398 9304 3662 9316
rect 3398 9096 3404 9304
rect 3612 9098 3662 9304
rect 3612 9096 3618 9098
rect -578 8532 -334 8538
rect -578 8312 -566 8532
rect -346 8312 -334 8532
rect 5664 8432 5752 8438
rect 5664 8368 5676 8432
rect 5740 8426 7858 8432
rect 5740 8374 7794 8426
rect 7846 8374 7858 8426
rect 5740 8368 7858 8374
rect 5664 8362 5752 8368
rect -578 8306 -334 8312
rect 3386 7884 3398 8110
rect 3618 7884 3630 8110
rect 3386 7878 3630 7884
rect 5254 7892 5330 7904
rect 7354 7892 7430 7898
rect 5254 7828 5260 7892
rect 5324 7886 5738 7892
rect 5324 7834 5674 7886
rect 5726 7834 5738 7886
rect 5324 7828 5738 7834
rect 7354 7828 7360 7892
rect 7424 7828 7430 7892
rect 5254 7816 5392 7828
rect 7354 7822 7430 7828
rect 5328 6646 5392 7816
rect 7360 6974 7424 7822
rect 7360 6910 8756 6974
rect 5328 6594 5334 6646
rect 5386 6594 5392 6646
rect 5328 6582 5392 6594
rect 7360 6646 7424 6910
rect 7360 6594 7366 6646
rect 7418 6594 7424 6646
rect 5670 6586 5746 6592
rect 5670 6522 5676 6586
rect 5740 6522 6452 6586
rect 7360 6582 7424 6594
rect 7764 6594 7852 6600
rect 7764 6530 7776 6594
rect 7840 6530 8980 6594
rect 7764 6524 7852 6530
rect 5670 6516 5746 6522
rect 5254 6298 5330 6304
rect 5254 6234 5260 6298
rect 5324 6292 7418 6298
rect 5324 6240 7354 6292
rect 7406 6240 7418 6292
rect 5324 6234 7418 6240
rect 5254 6228 5330 6234
rect 6408 5652 6472 6234
rect 6408 5588 6708 5652
rect 6772 5588 7432 5652
rect 5764 5280 5876 5292
rect 5764 5180 5770 5280
rect 5870 5204 6130 5280
rect 5870 5180 6036 5204
rect 5764 5168 5876 5180
rect 6030 5116 6036 5180
rect 6124 5116 6130 5204
rect 7368 5246 7432 5588
rect 7368 5194 7374 5246
rect 7426 5194 7432 5246
rect 7368 5182 7432 5194
rect 6030 5104 6130 5116
rect 5638 4898 5714 4904
rect 5638 4834 5644 4898
rect 5708 4892 6398 4898
rect 5708 4840 6334 4892
rect 6386 4840 6398 4892
rect 5708 4834 6398 4840
rect 5638 4828 5714 4834
rect 4960 4546 5056 4552
rect 4960 4474 4972 4546
rect 5044 4474 5056 4546
rect 4960 4468 5056 4474
rect 4972 2656 5044 4468
rect 4244 2584 5044 2656
rect 4094 1987 4167 1993
rect 4094 1908 4167 1914
rect 3034 1831 3124 1837
rect 3034 1825 3046 1831
rect 3034 1747 3040 1825
rect 3034 1741 3046 1747
rect 3124 1741 3130 1831
rect 3034 1735 3124 1741
rect 4244 1248 4316 2584
rect 5929 2250 5992 4834
rect 6054 4612 6130 4624
rect 8448 4612 8512 4618
rect 6054 4548 6060 4612
rect 6124 4606 8512 4612
rect 6124 4554 8454 4606
rect 8506 4554 8512 4606
rect 6124 4548 8512 4554
rect 6054 4536 6130 4548
rect 8448 4542 8512 4548
rect 8032 4334 8120 4340
rect 8032 4270 8044 4334
rect 8108 4328 8818 4334
rect 8108 4276 8754 4328
rect 8806 4276 8818 4328
rect 8108 4270 8818 4276
rect 8032 4264 8120 4270
rect 5929 2064 5992 2187
rect 8368 2282 8432 4270
rect 5728 2044 5986 2064
rect 5916 2006 5986 2044
rect 8368 2026 8432 2218
rect 5916 1955 5935 2006
rect 5916 1856 5986 1955
rect 8368 1974 8374 2026
rect 8426 1974 8432 2026
rect 8368 1956 8432 1974
rect 8368 1886 8432 1892
rect 5728 1768 5986 1856
rect -454 1242 4316 1248
rect -454 1182 -442 1242
rect -382 1182 4316 1242
rect -454 1176 4316 1182
rect 3478 1170 3550 1176
rect 3478 1110 3490 1170
rect 3478 1104 3550 1110
<< via1 >>
rect 6487 6906 6585 6912
rect 6487 6820 6493 6906
rect 6493 6820 6579 6906
rect 6579 6820 6585 6906
rect 6487 6814 6585 6820
rect 6708 5588 6772 5652
rect 3046 1825 3124 1831
rect 3046 1747 3118 1825
rect 3118 1747 3124 1825
rect 3046 1741 3124 1747
rect 5929 2187 5992 2250
rect 8368 2218 8432 2282
rect 4529 1975 4590 1981
rect 4529 1926 4535 1975
rect 4535 1926 4584 1975
rect 4584 1926 4590 1975
rect 4529 1920 4590 1926
rect 6708 2006 6772 2012
rect 6708 1954 6714 2006
rect 6714 1954 6766 2006
rect 6766 1954 6772 2006
rect 6708 1948 6772 1954
rect 8368 1950 8432 1956
rect 8368 1898 8374 1950
rect 8374 1898 8426 1950
rect 8426 1898 8432 1950
rect 8368 1892 8432 1898
<< metal2 >>
rect 6493 6453 6579 6814
rect 5923 2187 5929 2250
rect 5992 2187 5998 2250
rect 4522 2120 4590 2122
rect 5929 2120 5992 2187
rect 6494 2120 6579 6453
rect 8362 2218 8368 2282
rect 8432 2218 8438 2282
rect 8368 2120 8432 2218
rect 4522 1981 6708 2120
rect 4590 1948 6708 1981
rect 6772 1956 9234 2120
rect 6772 1948 8368 1956
rect 4590 1920 8368 1948
rect 4522 1892 8368 1920
rect 8432 1892 9234 1956
rect 3046 1831 3124 1837
rect 4522 1825 9234 1892
rect 3124 1747 9234 1825
rect 3046 1735 3124 1741
rect 4522 1518 9234 1747
<< metal3 >>
rect 4824 2090 5144 2091
rect 4824 1772 4825 2090
rect 5143 1772 5144 2090
rect 4824 1771 5144 1772
<< metal5 >>
rect 4800 2091 5168 2115
rect 4800 1771 4824 2091
rect 5144 1771 5168 2091
rect 4800 1747 5168 1771
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_0 ~/aicex/ip/cnr_gr00_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 4684 0 1 5824
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_1
timestamp 1695852000
transform 1 0 6784 0 1 5824
box -184 -124 1528 1016
use CNRATR_NCH_8C4F0  CNRATR_NCH_8C4F0_0 ~/aicex/ip/cnr_gr00_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 4684 0 1 4424
box -184 -124 1912 1016
use CNRATR_NCH_8C12F0  CNRATR_NCH_8C12F0_0 ~/aicex/ip/cnr_gr00_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 7084 0 1 3284
box -184 -124 1912 2168
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_0 ~/aicex/ip/cnr_gr00_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 6784 0 1 7124
box -184 -124 1528 1592
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_1
timestamp 1695852000
transform 1 0 4684 0 1 7124
box -184 -124 1528 1592
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712309819
transform 0 -1 3092 1 0 428
box 0 0 8720 4236
<< labels >>
flabel locali 3612 9100 8200 9300 0 FreeSans 1600 0 0 0 VDD_1V8
port 1 nsew
flabel metal1 7840 6530 8980 6594 0 FreeSans 1600 0 0 0 VIN
port 3 nsew
flabel metal1 5740 6522 6452 6586 0 FreeSans 1600 0 0 0 VIP
port 4 nsew
flabel metal1 7360 6910 8756 6974 0 FreeSans 1600 0 0 0 OPAMP_VOUT
port 5 nsew
flabel metal2 4522 1518 9234 1890 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
<< end >>

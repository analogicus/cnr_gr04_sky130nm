*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_GR04_T2I_S_lpe.spi
#else
.include ../../../work/xsch/CNR_GR04_T2I_S.spice
.include ../../../design/time-to-digital/SPICE/top.cir
#endif
.include ../../../design/time-to-digital/HDL/runs/RUN_2024-04-12_12-12-37/final/spice/top.spice

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15
.option TEMP=27

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param AVDD = {vdda}

*Controller CLK
.param CLK_FREQ = 20MEG
.param PERIOD = 1/CLK_FREQ
.param HALF_PERIOD = PERIOD/2

*Simulation Control
.param SIM_STEP = 1n
.param SIM_START = 1n
.param SIM_STOP = 100000000000*PERIOD


*Inputs
.param RESET_START = 2*PERIOD
.param START = 4*PERIOD
.param DATA_HALF_PERIOD = 10*PERIOD
.param DATA_PERIOD = 20*PERIOD

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  dc 1.8

*VRESET RESET 0 pulse 0 1.8 0 0 0 50ns 2000ns

R_reset RESET temp_reset 0

VCLK    CLK     VSS   PULSE(0 1.8 0           0 0 HALF_PERIOD PERIOD)
VRST    RST     VSS   PULSE(0 1.8 RESET_START 0 0 PERIOD SIM_STOP)
VSTART  START   VSS   PULSE(0 1.8 START       0 0 PERIOD SIM_STOP)
*VDATA   data_in VSS   PULSE(0 1.8 0          0 0 DATA_HALF_PERIOD DATA_PERIOD)




*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
*XU1 CLK RST COMPERATOR START ready running temp_reset d7 d6 d5 d4 d3 d2 d1 d0 top_verilog

XU2 VSS VDD_1V8 CLK d0 d1 d2 d3 d4 d5 d6 COMPERATOR ready RST running START temp_reset top


R0 d0 VDD_1V8 1k
R1 d1 VDD_1V8 1k
R2 d2 VDD_1V8 1k
R3 d3 VDD_1V8 1k
R4 d4 VDD_1V8 1k
R5 d5 VDD_1V8 1k
R6 d6 VDD_1V8 1k
R7 d7 VDD_1V8 1k

R_Running running VDD_1V8 1k


*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------

.save V(CLK) V(RST) V(COMPERATOR) V(START)
.save V(temp_reset) V(ready) V(running)
.save V(d7) V(d6) V(d5) V(d4) V(d3) V(d2) V(d1) V(d0)
.save V(VDD) -I(VDD)
.save all
*----------------------------------------------------------------

* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save ${VPORTS} 
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 1 1 1 100p 20u 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else

*tran 1n 400u 1p
tran 1n 20u 0
    
*dc TEMP -40 125 1
write

*plot V(CLK_OUT)
*Controlller input
plot V(RST) V(START) V(COMPERATOR)

*Controller output
*plot V(ready) V(running) V(temp_reset) 
*plot V(running) V(COMPERATOR)
*plot V(d7) V(d6) V(d5) V(d4) V(d3) V(d2) V(d1) V(d0)
quit
#endif
.endc
.end

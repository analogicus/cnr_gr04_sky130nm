magic
tech sky130B
magscale 1 2
timestamp 1713440215
<< metal4 >>
rect -7447 2039 -2749 2080
rect -7447 -2039 -3005 2039
rect -2769 -2039 -2749 2039
rect -7447 -2080 -2749 -2039
rect -2349 2039 2349 2080
rect -2349 -2039 2093 2039
rect 2329 -2039 2349 2039
rect -2349 -2080 2349 -2039
rect 2749 2039 7447 2080
rect 2749 -2039 7191 2039
rect 7427 -2039 7447 2039
rect 2749 -2080 7447 -2039
<< via4 >>
rect -3005 -2039 -2769 2039
rect 2093 -2039 2329 2039
rect 7191 -2039 7427 2039
<< mimcap2 >>
rect -7367 1960 -3367 2000
rect -7367 -1960 -7327 1960
rect -3407 -1960 -3367 1960
rect -7367 -2000 -3367 -1960
rect -2269 1960 1731 2000
rect -2269 -1960 -2229 1960
rect 1691 -1960 1731 1960
rect -2269 -2000 1731 -1960
rect 2829 1960 6829 2000
rect 2829 -1960 2869 1960
rect 6789 -1960 6829 1960
rect 2829 -2000 6829 -1960
<< mimcap2contact >>
rect -7327 -1960 -3407 1960
rect -2229 -1960 1691 1960
rect 2869 -1960 6789 1960
<< metal5 >>
rect -3047 2039 -2727 2081
rect -7351 1960 -3383 1984
rect -7351 -1960 -7327 1960
rect -3407 -1960 -3383 1960
rect -7351 -1984 -3383 -1960
rect -3047 -2039 -3005 2039
rect -2769 -2039 -2727 2039
rect 2051 2039 2371 2081
rect -2253 1960 1715 1984
rect -2253 -1960 -2229 1960
rect 1691 -1960 1715 1960
rect -2253 -1984 1715 -1960
rect -3047 -2081 -2727 -2039
rect 2051 -2039 2093 2039
rect 2329 -2039 2371 2039
rect 7149 2039 7469 2081
rect 2845 1960 6813 1984
rect 2845 -1960 2869 1960
rect 6789 -1960 6813 1960
rect 2845 -1984 6813 -1960
rect 2051 -2081 2371 -2039
rect 7149 -2039 7191 2039
rect 7427 -2039 7469 2039
rect 7149 -2081 7469 -2039
<< properties >>
string FIXED_BBOX 2749 -2080 6909 2080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20.0 l 20.0 val 815.2 carea 2.00 cperi 0.19 nx 3 ny 1 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1713508964
<< error_p >>
rect 23780 13822 23786 13824
rect 23857 13822 23863 13824
rect 23780 13819 23794 13822
rect 23849 13819 23863 13822
rect 23780 13818 23786 13819
rect 23857 13818 23863 13819
rect 23774 13813 23869 13818
rect 23774 13812 23785 13813
rect 23638 13667 23694 13811
rect 23776 13804 23785 13812
rect 23858 13812 23869 13813
rect 23858 13804 23867 13812
rect 23780 13749 23785 13804
rect 23776 13741 23785 13749
rect 23774 13740 23785 13741
rect 23858 13741 23867 13749
rect 23858 13740 23869 13741
rect 23774 13735 23869 13740
rect 23780 13734 23786 13735
rect 23857 13734 23863 13735
rect 23780 13731 23794 13734
rect 23849 13731 23863 13734
rect 23780 13729 23786 13731
rect 23857 13729 23863 13731
rect 23638 13617 23982 13667
rect 23638 13593 23694 13617
rect 23602 13557 24042 13587
rect 23318 13273 23694 13491
rect 27506 13380 27512 13392
rect 27588 13380 27594 13392
rect 27518 13368 27530 13374
rect 27570 13368 27582 13374
rect 27570 12802 27582 12808
rect 27588 12784 27594 12796
rect 27588 12732 27594 12744
rect 27570 12720 27582 12726
rect 27934 12230 27946 12236
rect 27986 12230 27998 12236
rect 27922 12212 27928 12224
rect 28004 12212 28010 12224
rect 26963 11990 27038 11993
rect 28190 11990 28253 11993
rect 26963 11956 27072 11959
rect 28156 11956 28253 11959
rect 41620 10896 41626 10908
rect 41858 10896 41864 10908
rect 41632 10884 41644 10890
rect 41840 10884 41852 10890
rect 47557 10854 47563 10866
rect 47661 10854 47667 10866
rect 47569 10842 47581 10848
rect 47643 10842 47655 10848
rect 46930 10771 46942 10777
rect 46918 10753 46924 10765
rect 46918 10701 46924 10713
rect 46930 10689 46942 10695
rect 530 10498 536 10510
rect 768 10498 774 10510
rect 542 10486 554 10492
rect 750 10486 762 10492
rect 6467 10456 6473 10468
rect 6571 10456 6577 10468
rect 6479 10444 6491 10450
rect 6553 10444 6565 10450
rect 20129 10437 20135 10449
rect 20233 10437 20239 10449
rect 20141 10425 20153 10431
rect 20215 10425 20227 10431
rect 5840 10373 5852 10379
rect 5828 10355 5834 10367
rect 5828 10303 5834 10315
rect 5840 10291 5852 10297
rect 47554 8994 47572 9000
rect 47634 8994 47652 9000
rect 47548 8976 47554 8994
rect 47652 8976 47658 8994
rect 47548 8896 47554 8914
rect 47652 8896 47658 8914
rect 47554 8890 47572 8896
rect 47634 8890 47652 8896
rect 46502 8710 46508 8722
rect 46584 8710 46590 8722
rect 48924 8712 48942 8718
rect 48982 8712 49000 8718
rect 46514 8698 46526 8704
rect 46566 8698 46578 8704
rect 48918 8694 48924 8712
rect 49000 8694 49006 8712
rect 48918 8636 48924 8654
rect 49000 8636 49006 8654
rect 48924 8630 48942 8636
rect 48982 8630 49000 8636
rect 6464 8596 6482 8602
rect 6544 8596 6562 8602
rect 6458 8578 6464 8596
rect 6562 8578 6568 8596
rect 6458 8498 6464 8516
rect 6562 8498 6568 8516
rect 6464 8492 6482 8498
rect 6544 8492 6562 8498
rect 12717 8478 12720 8484
rect 17080 8478 17092 8484
rect 17288 8478 17300 8484
rect 12729 8460 12732 8472
rect 17068 8460 17074 8472
rect 17306 8460 17312 8472
rect 5412 8312 5418 8324
rect 5494 8312 5500 8324
rect 7840 8314 7852 8320
rect 5424 8300 5436 8306
rect 5476 8300 5488 8306
rect 7828 8296 7834 8308
rect 7828 8244 7834 8256
rect 12729 8252 12732 8264
rect 15388 8252 15394 8264
rect 15626 8252 15632 8264
rect 18288 8252 18294 8264
rect 18526 8252 18532 8264
rect 12708 8240 12720 8246
rect 15400 8240 15412 8246
rect 15608 8240 15620 8246
rect 18300 8240 18312 8246
rect 18508 8240 18520 8246
rect 7840 8232 7852 8238
rect 9720 8001 9721 8007
rect 9708 7983 9714 7995
rect 9720 7934 9782 7960
rect 9682 7896 9694 7922
rect 9760 7896 9794 7922
rect 9660 7388 9694 7398
rect 9760 7388 9782 7398
rect 9681 7350 9744 7360
rect 9669 7301 9675 7313
rect 9750 7301 9756 7313
rect 9681 7289 9683 7295
rect 9742 7289 9744 7295
rect 47302 7139 47308 7151
rect 47384 7139 47390 7151
rect 47314 7127 47326 7133
rect 47366 7127 47378 7133
rect 6212 6741 6218 6753
rect 6294 6741 6300 6753
rect 6224 6729 6236 6735
rect 6276 6729 6288 6735
rect 9683 6634 9742 6635
rect 9660 6600 9742 6634
rect 9760 6600 9780 6634
rect 9683 6576 9742 6600
rect 47302 5667 47308 5679
rect 47384 5667 47390 5679
rect 47314 5655 47326 5661
rect 47366 5655 47378 5661
rect 9683 5346 9742 5349
rect 9660 5312 9742 5346
rect 9760 5312 9780 5346
rect 9683 5290 9742 5312
rect 6212 5269 6218 5281
rect 6294 5269 6300 5281
rect 6224 5257 6236 5263
rect 6276 5257 6288 5263
rect 46758 4898 46770 4904
rect 46776 4880 46782 4892
rect 46776 4828 46782 4840
rect 46758 4816 46770 4822
rect 5668 4500 5680 4506
rect 5686 4482 5692 4494
rect 5686 4430 5692 4442
rect 5668 4418 5680 4424
rect 13465 4280 13471 4292
rect 13631 4280 13637 4292
rect 13477 4268 13489 4274
rect 13613 4268 13625 4274
rect 13165 3910 13175 3929
rect 14450 3910 14463 3929
rect 15740 3910 15751 3929
rect 17026 3910 17039 3929
rect 18318 3910 18327 3929
rect 19606 3910 19615 3929
rect 20891 3910 20903 3929
rect 13250 3897 13262 3903
rect 20976 3897 20988 3903
rect 13165 3810 13175 3844
rect 13203 3830 13213 3891
rect 13268 3890 13274 3891
rect 13268 3830 13274 3831
rect 13250 3818 13262 3824
rect 14450 3810 14463 3844
rect 14488 3831 14501 3891
rect 15740 3810 15751 3844
rect 15778 3832 15789 3891
rect 17026 3810 17039 3844
rect 17064 3832 17077 3891
rect 18318 3810 18327 3844
rect 18356 3832 18365 3891
rect 19606 3810 19615 3844
rect 19644 3832 19653 3891
rect 20891 3810 20903 3844
rect 20929 3832 20941 3891
rect 20994 3879 21000 3891
rect 20994 3832 21000 3844
rect 20976 3820 20988 3826
rect 25812 723 25838 747
rect 26216 668 26452 676
rect 26096 627 26472 652
rect 26132 597 26158 616
rect 26132 595 26163 597
rect 26473 595 26479 597
rect 26132 592 26171 595
rect 26465 592 26479 595
rect 26156 591 26480 592
rect 26151 585 26485 591
rect 26153 577 26483 585
rect 26156 547 26480 577
rect 26153 275 26162 283
rect 26151 274 26162 275
rect 26474 275 26483 283
rect 26474 274 26485 275
rect 26151 269 26157 274
rect 26162 269 26171 274
rect 26157 265 26171 269
rect 26465 269 26474 274
rect 26479 269 26485 274
rect 26465 265 26479 269
rect 26157 263 26163 265
rect 26473 263 26479 265
<< error_s >>
rect 10485 10380 10491 10392
rect 10589 10380 10595 10392
rect 10497 10368 10509 10374
rect 10571 10368 10583 10374
rect 9840 10306 9852 10312
rect 9828 10288 9834 10300
rect 9828 10236 9834 10248
rect 9840 10224 9852 10230
rect 9683 4063 9742 4088
rect 9660 4029 9742 4063
rect 9660 4024 9694 4029
rect 9760 4024 9780 4058
<< locali >>
rect 9206 2614 10394 2914
<< metal1 >>
rect 9734 11014 11860 11314
use CNR_GR04_T2I_S  CNR_GR04_T2I_S_0
timestamp 1713464657
transform 1 0 -36 0 1 2614
box 0 -2598 49502 12158
<< labels >>
flabel locali 9416 2614 9716 2914 0 FreeSans 1600 0 0 0 VSS
port 3 nsew
<< end >>

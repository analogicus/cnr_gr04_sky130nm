magic
tech sky130B
magscale 1 2
timestamp 1713447325
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__pfet_01v8_GYUYCA  XM1
timestamp 0
transform 1 0 280 0 1 958
box 0 0 1 1
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 D
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 G
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 S
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 B
port 3 nsew
<< end >>

magic
tech sky130B
magscale 1 2
timestamp 1712903178
<< error_s >>
rect 754 1847 760 1853
rect 825 1847 831 1853
rect 748 1841 754 1847
rect 831 1841 837 1847
rect 2972 1846 2990 1852
rect 3030 1846 3048 1852
rect 2966 1828 2972 1846
rect 3048 1828 3054 1846
rect 748 1770 754 1776
rect 831 1770 837 1776
rect 2966 1770 2972 1788
rect 3048 1770 3054 1788
rect 754 1764 760 1770
rect 825 1764 831 1770
rect 2972 1764 2990 1770
rect 3030 1764 3048 1770
rect 2126 -641 2135 -632
rect 2182 -641 2191 -632
rect 2550 -637 2559 -633
rect 2605 -637 2614 -633
rect 2117 -642 2126 -641
rect 2191 -642 2200 -641
rect 2545 -642 2619 -637
rect 2117 -650 2120 -642
rect 2196 -650 2200 -642
rect 2541 -651 2544 -642
rect 2117 -706 2120 -697
rect 2196 -706 2200 -697
rect 2541 -706 2544 -697
rect 2545 -706 2550 -642
rect 2620 -651 2623 -642
rect 2620 -706 2623 -697
rect 2126 -715 2135 -706
rect 2182 -715 2191 -706
rect 2545 -711 2619 -706
rect 2550 -715 2559 -711
rect 2605 -715 2614 -711
rect 965 -811 977 -805
rect 987 -811 999 -805
rect 953 -829 959 -817
rect 1005 -818 1011 -817
rect 953 -851 959 -839
rect 1005 -851 1011 -850
rect 965 -863 977 -857
rect 987 -863 999 -857
rect 1428 -2936 1482 -2920
rect 1456 -2964 1482 -2948
rect 1237 -3259 1249 -3253
rect 1259 -3259 1271 -3253
rect 1225 -3277 1231 -3265
rect 1277 -3266 1283 -3265
rect 1225 -3299 1231 -3287
rect 1277 -3299 1283 -3298
rect 1237 -3311 1249 -3305
rect 1259 -3311 1271 -3305
rect -4558 -3436 -4524 -3418
rect -4530 -3478 -4524 -3460
rect 3701 -3501 3713 -3495
rect 3723 -3501 3735 -3495
rect 3854 -3498 3860 -3492
rect 3900 -3498 3906 -3492
rect 3848 -3504 3854 -3498
rect 3906 -3504 3912 -3498
rect 3689 -3519 3695 -3507
rect 3741 -3508 3747 -3507
rect 3689 -3541 3695 -3529
rect 3741 -3541 3747 -3540
rect 3701 -3553 3713 -3547
rect 3723 -3553 3735 -3547
rect 3848 -3550 3854 -3544
rect 3906 -3550 3912 -3544
rect 3854 -3556 3860 -3550
rect 3900 -3556 3906 -3550
rect 374 -3596 386 -3590
rect 434 -3596 446 -3590
rect 362 -3614 368 -3602
rect 452 -3614 458 -3602
rect -4548 -3766 -4514 -3748
rect -4520 -3808 -4514 -3790
rect 2128 -5280 2134 -5274
rect 2182 -5280 2188 -5274
rect 2122 -5286 2128 -5280
rect 2188 -5286 2194 -5280
rect 2122 -5340 2128 -5336
rect 2188 -5340 2194 -5336
rect 2128 -5346 2134 -5340
rect 2182 -5346 2188 -5340
<< locali >>
rect 958 2477 984 2496
rect 958 2424 984 2443
rect 3640 -700 3642 -648
<< viali >>
rect 951 2443 985 2477
rect 1513 2443 1547 2477
rect 3169 2445 3203 2479
rect 3731 2445 3765 2479
rect -1174 1862 -954 2082
rect 760 1776 825 1841
rect 951 1791 985 1825
rect 1195 1791 1229 1825
rect 2978 1776 3042 1840
rect 1176 1272 1240 1336
rect 3398 1278 3450 1330
rect 766 -506 819 -453
rect 2984 -500 3036 -448
rect 1574 -706 1638 -642
rect 3642 -700 3692 -648
rect 965 -851 999 -817
rect 2801 -851 2835 -817
rect -4574 -2488 -4522 -2436
rect 2878 -2620 2918 -2580
rect 1237 -2937 1271 -2903
rect 1462 -3024 1526 -2960
rect 3922 -3018 3974 -2966
rect 1237 -3299 1271 -3265
rect 1727 -3299 1761 -3265
rect 3701 -3541 3735 -3507
rect 4189 -3541 4223 -3507
rect 374 -3674 446 -3602
rect -1094 -5082 -1034 -5022
<< metal1 >>
rect -1272 3018 3776 3336
rect -1174 2088 -954 3018
rect 945 2477 991 2489
rect 945 2443 951 2477
rect 985 2476 991 2477
rect 1198 2476 1230 3018
rect 1501 2477 1559 2483
rect 1501 2476 1513 2477
rect 985 2444 1513 2476
rect 985 2443 991 2444
rect 945 2431 991 2443
rect 1501 2443 1513 2444
rect 1547 2443 1559 2477
rect 1501 2437 1559 2443
rect 3163 2479 3209 2491
rect 3163 2445 3169 2479
rect 3203 2478 3209 2479
rect 3408 2478 3440 3018
rect 3719 2479 3777 2485
rect 3719 2478 3731 2479
rect 3203 2446 3731 2478
rect 3203 2445 3209 2446
rect 3163 2433 3209 2445
rect 3719 2445 3731 2446
rect 3765 2445 3777 2479
rect 3719 2439 3777 2445
rect -1186 2082 -942 2088
rect -1186 1862 -1174 2082
rect -954 1862 -942 2082
rect -1186 1856 -942 1862
rect 754 1847 831 1853
rect 945 1825 991 1837
rect 945 1791 951 1825
rect 985 1824 991 1825
rect 1183 1825 1241 1831
rect 1183 1824 1195 1825
rect 985 1792 1195 1824
rect 985 1791 991 1792
rect 945 1779 991 1791
rect 1183 1791 1195 1792
rect 1229 1791 1241 1825
rect 1183 1785 1241 1791
rect 754 1764 831 1770
rect 1170 1336 1246 1348
rect 1170 1272 1176 1336
rect 1240 1330 3462 1336
rect 1240 1278 3398 1330
rect 3450 1278 3462 1330
rect 1240 1272 3462 1278
rect 1170 1260 1246 1272
rect 754 -512 760 -447
rect 825 -512 831 -447
rect 2972 -506 2978 -442
rect 3042 -506 3048 -442
rect 1568 -642 1644 -630
rect 2126 -642 2190 -636
rect 2550 -642 2614 -636
rect 1568 -706 1574 -642
rect 1638 -706 2126 -642
rect 2190 -706 2550 -642
rect 2614 -648 3704 -642
rect 2614 -700 3642 -648
rect 3692 -700 3704 -648
rect 2614 -706 3704 -700
rect 1568 -718 1644 -706
rect 2126 -712 2190 -706
rect 2550 -712 2614 -706
rect 1928 -808 1980 -802
rect 959 -817 1005 -811
rect 959 -851 965 -817
rect 999 -818 1005 -817
rect 999 -850 1928 -818
rect 999 -851 1005 -850
rect 959 -857 1005 -851
rect 2795 -817 2841 -805
rect 2795 -818 2801 -817
rect 1980 -850 2801 -818
rect 1928 -866 1980 -860
rect 2795 -851 2801 -850
rect 2835 -851 2841 -817
rect 2795 -863 2841 -851
rect -4586 -2436 2218 -2430
rect -4586 -2488 -4574 -2436
rect -4522 -2488 2218 -2436
rect -4586 -2494 2218 -2488
rect 1231 -2903 1277 -2891
rect 1231 -2937 1237 -2903
rect 1271 -2904 1277 -2903
rect 1271 -2936 1514 -2904
rect 1271 -2937 1277 -2936
rect 1231 -2949 1277 -2937
rect 1482 -2948 1514 -2936
rect 1456 -2960 1532 -2948
rect 2154 -2960 2218 -2494
rect 2866 -2626 2872 -2574
rect 2924 -2626 2930 -2574
rect 3916 -2960 3980 -2954
rect 1456 -3024 1462 -2960
rect 1526 -2966 3980 -2960
rect 1526 -3018 3922 -2966
rect 3974 -3018 3980 -2966
rect 1526 -3024 3980 -3018
rect 1456 -3036 1532 -3024
rect 3916 -3030 3980 -3024
rect 1384 -3256 1436 -3250
rect 1231 -3265 1277 -3259
rect 1231 -3299 1237 -3265
rect 1271 -3266 1277 -3265
rect 1271 -3298 1384 -3266
rect 1271 -3299 1277 -3298
rect 1231 -3305 1277 -3299
rect 1715 -3265 1773 -3259
rect 1715 -3266 1727 -3265
rect 1436 -3298 1727 -3266
rect 1384 -3314 1436 -3308
rect -4582 -3436 -4530 -3430
rect -4582 -3494 -4530 -3488
rect 368 -3602 452 -3596
rect 368 -3674 374 -3602
rect 446 -3674 452 -3602
rect 368 -3680 452 -3674
rect -4572 -3766 -4520 -3760
rect -4572 -3824 -4520 -3818
rect 374 -5016 446 -3680
rect -1106 -5022 446 -5016
rect -1106 -5082 -1094 -5022
rect -1034 -5082 446 -5022
rect -1106 -5088 446 -5082
rect 1608 -5304 1640 -3298
rect 1715 -3299 1727 -3298
rect 1761 -3299 1773 -3265
rect 1715 -3305 1773 -3299
rect 3695 -3507 3741 -3501
rect 3695 -3541 3701 -3507
rect 3735 -3508 3741 -3507
rect 3735 -3540 3854 -3508
rect 3735 -3541 3741 -3540
rect 3695 -3547 3741 -3541
rect 4096 -3508 4128 -3504
rect 4177 -3507 4235 -3501
rect 4177 -3508 4189 -3507
rect 3906 -3540 4189 -3508
rect 1608 -5336 2128 -5304
rect 4096 -5304 4128 -3540
rect 4177 -3541 4189 -3540
rect 4223 -3541 4235 -3507
rect 4177 -3547 4235 -3541
rect 2188 -5336 4128 -5304
<< via1 >>
rect 754 1841 831 1847
rect 754 1776 760 1841
rect 760 1776 825 1841
rect 825 1776 831 1841
rect 2972 1840 3048 1846
rect 754 1770 831 1776
rect 2972 1776 2978 1840
rect 2978 1776 3042 1840
rect 3042 1776 3048 1840
rect 2972 1770 3048 1776
rect 760 -453 825 -447
rect 760 -506 766 -453
rect 766 -506 819 -453
rect 819 -506 825 -453
rect 760 -512 825 -506
rect 2978 -448 3042 -442
rect 2978 -500 2984 -448
rect 2984 -500 3036 -448
rect 3036 -500 3042 -448
rect 2978 -506 3042 -500
rect 2126 -706 2190 -642
rect 2550 -706 2614 -642
rect 1928 -860 1980 -808
rect 2872 -2580 2924 -2574
rect 2872 -2620 2878 -2580
rect 2878 -2620 2918 -2580
rect 2918 -2620 2924 -2580
rect 2872 -2626 2924 -2620
rect 1384 -3308 1436 -3256
rect -4582 -3488 -4530 -3436
rect -4572 -3818 -4520 -3766
rect 3854 -3550 3906 -3498
rect 2128 -5340 2188 -5280
<< metal2 >>
rect 760 -447 825 1770
rect 2978 -442 3042 1770
rect 2978 -512 3042 -506
rect 760 -518 825 -512
rect 2120 -706 2126 -642
rect 2191 -706 2196 -642
rect 2544 -706 2550 -642
rect 2614 -706 2620 -642
rect 1922 -860 1928 -808
rect 1980 -860 1986 -808
rect 1938 -1554 1970 -860
rect 1938 -1586 2914 -1554
rect 2882 -2568 2914 -1586
rect 2872 -2574 2924 -2568
rect 2872 -2632 2924 -2626
rect 1378 -3308 1384 -3256
rect 1436 -3308 1442 -3256
rect -4588 -3488 -4582 -3436
rect -4530 -3446 -4524 -3436
rect -4530 -3488 -4524 -3478
rect -4578 -3818 -4572 -3766
rect -4520 -3776 -4514 -3766
rect -4520 -3818 -4514 -3808
rect 2121 -5338 2128 -5282
rect 2188 -5338 2195 -5282
<< via2 >>
rect 2126 -642 2191 -641
rect 2126 -706 2190 -642
rect 2190 -706 2191 -642
rect 2550 -706 2614 -642
rect 2130 -5338 2186 -5282
<< metal3 >>
rect 2121 -641 2196 -636
rect 2121 -706 2126 -641
rect 2191 -706 2196 -641
rect 2121 -711 2196 -706
rect 2545 -642 2619 -637
rect 2545 -706 2550 -642
rect 2614 -706 2619 -642
rect 2545 -711 2619 -706
rect 2126 -1182 2191 -711
rect 2128 -5277 2188 -1182
rect 2125 -5282 2191 -5277
rect 2125 -5338 2130 -5282
rect 2186 -5338 2191 -5282
rect 2125 -5343 2191 -5338
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 2392 0 1 -1284
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_1
timestamp 1695852000
transform 1 0 198 0 1 -1284
box -184 -124 1528 1016
use CNRATR_NCH_8C4F0  CNRATR_NCH_8C4F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 86 0 1 -3724
box -184 -124 1912 1016
use CNRATR_NCH_8C12F0  CNRATR_NCH_8C12F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 2550 0 1 -4546
box -184 -124 1912 2168
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 2402 0 1 1078
box -184 -124 1528 1592
use CNRATR_PCH_4C8F0  CNRATR_PCH_4C8F0_1
timestamp 1695852000
transform 1 0 184 0 1 1078
box -184 -124 1528 1592
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/sun_tr_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712309819
transform 0 1 -4612 -1 0 2698
box 0 0 8720 4236
<< labels >>
flabel metal1 -1272 3018 3776 3336 0 FreeSans 1600 0 0 0 VDD_1V8
port 6 nsew
flabel space 3384 -586 3448 -514 0 FreeSans 160 0 0 0 VIN
port 3 nsew
flabel metal1 1640 -706 3642 -642 0 FreeSans 160 0 0 0 VSS
port 7 nsew
flabel metal1 1608 -5336 4128 -5304 0 FreeSans 160 0 0 0 VSS
port 8 nsew
flabel space 1188 -586 1252 -514 0 FreeSans 160 0 0 0 VIP
port 9 nsew
flabel metal2 2978 -442 3042 1770 0 FreeSans 160 0 0 0 OPAMP_VOUT
port 10 nsew
<< end >>

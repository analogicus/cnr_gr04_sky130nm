magic
tech sky130B
magscale 1 2
timestamp 1713473354
<< error_s >>
rect 775 418 812 421
rect 809 393 812 399
rect 840 393 843 399
rect 803 390 812 393
rect 797 375 803 387
rect 849 375 855 387
rect 797 353 803 365
rect 849 353 855 365
rect 809 341 821 347
rect 831 341 843 347
rect 1580 -98 1584 639
rect 6077 321 6089 327
rect 6099 321 6111 327
rect 6065 303 6071 315
rect 6117 314 6123 315
rect 6065 281 6071 293
rect 6117 281 6123 282
rect 6077 269 6089 275
rect 6099 269 6111 275
rect 4608 -374 4617 -367
rect 4659 -374 4668 -367
rect 4608 -376 4612 -374
rect 4664 -376 4668 -374
rect 4599 -385 4608 -376
rect 4668 -385 4677 -376
rect 1512 -400 1521 -391
rect 1563 -400 1572 -391
rect 1503 -404 1512 -400
rect 1572 -404 1581 -400
rect 1503 -409 1510 -404
rect 1574 -409 1581 -404
rect 7962 -404 7971 -397
rect 8013 -404 8022 -397
rect 7962 -406 7966 -404
rect 8018 -406 8022 -404
rect 7953 -415 7962 -406
rect 8022 -415 8031 -406
rect 4599 -436 4608 -427
rect 4668 -436 4677 -427
rect 4608 -438 4612 -436
rect 4664 -438 4668 -436
rect 4608 -445 4617 -438
rect 4659 -445 4668 -438
rect 1503 -456 1510 -451
rect 1574 -456 1581 -451
rect 1503 -460 1512 -456
rect 1572 -460 1581 -456
rect 1512 -469 1521 -460
rect 1563 -469 1572 -460
rect 7953 -466 7962 -457
rect 8022 -466 8031 -457
rect 7962 -468 7966 -466
rect 8018 -468 8022 -466
rect 7962 -475 7971 -468
rect 8013 -475 8022 -468
rect 9258 -938 9267 -935
rect 9473 -938 9482 -935
rect 9252 -944 9488 -938
rect 9249 -953 9491 -944
rect 9252 -962 9488 -953
rect 636 -1068 876 -1060
rect 1428 -1068 1668 -1060
rect 7130 -1079 7370 -1056
rect 7922 -1079 8162 -1056
rect 664 -1096 848 -1088
rect 1456 -1096 1640 -1088
rect 3792 -1110 4032 -1084
rect 4584 -1110 4824 -1084
rect 7158 -1107 7342 -1084
rect 7950 -1107 8134 -1084
rect 3820 -1138 4004 -1112
rect 4612 -1138 4796 -1112
rect 9252 -1150 9276 -962
rect 9464 -1150 9488 -962
rect 9252 -1159 9488 -1150
rect 9249 -1168 9491 -1159
rect 9252 -1174 9488 -1168
rect 9258 -1177 9267 -1174
rect 9473 -1177 9482 -1174
rect 7122 -1514 9671 -1357
rect 2955 -1611 3137 -1575
rect 2955 -1713 2991 -1611
rect 3101 -1713 3137 -1611
rect 7122 -1677 7158 -1514
rect 7442 -1635 9671 -1514
rect 7469 -1677 8477 -1659
rect 2955 -1749 3137 -1713
rect 670 -2173 694 -1855
rect 824 -1951 833 -1947
rect 875 -1951 884 -1947
rect 819 -1956 889 -1951
rect 815 -1965 818 -1956
rect 815 -2016 818 -2007
rect 819 -2016 824 -1956
rect 890 -1965 893 -1956
rect 890 -2016 893 -2007
rect 819 -2027 889 -2016
rect 1014 -2173 1038 -1855
rect 2238 -2156 2246 -2078
rect 2558 -2174 2582 -1758
rect 4467 -2087 4491 -1807
rect 4613 -1862 4619 -1860
rect 4682 -1862 4688 -1860
rect 4613 -1866 4627 -1862
rect 4674 -1866 4688 -1862
rect 4607 -1871 4694 -1866
rect 4607 -1872 4618 -1871
rect 4688 -1872 4694 -1871
rect 4609 -1880 4612 -1872
rect 4609 -1935 4612 -1927
rect 4613 -1935 4618 -1872
rect 4689 -1880 4692 -1872
rect 4689 -1935 4692 -1927
rect 4607 -1936 4618 -1935
rect 4688 -1936 4694 -1935
rect 4607 -1941 4694 -1936
rect 4613 -1945 4627 -1941
rect 4674 -1945 4688 -1941
rect 4613 -1947 4619 -1945
rect 4682 -1947 4688 -1945
rect 4811 -2087 4835 -1807
rect 6192 -1854 6216 -1710
rect 7442 -1795 7478 -1677
rect 7158 -1798 7478 -1795
rect 350 -2493 694 -2175
rect 1014 -2493 1358 -2175
rect 1918 -2476 1926 -2175
rect 4147 -2407 4491 -2127
rect 4811 -2407 5155 -2127
rect 5552 -2458 5560 -2127
rect 5872 -2138 5880 -2030
rect 6192 -2174 6216 -1979
rect 7789 -1997 8157 -1979
rect 9393 -2018 9671 -1635
rect 7813 -2099 8133 -2097
rect 6894 -2118 7762 -2115
rect 7922 -2128 8024 -2112
rect 7932 -2133 8024 -2128
rect 7932 -2134 7943 -2133
rect 8003 -2134 8024 -2133
rect 7934 -2139 7937 -2134
rect 7938 -2139 7943 -2134
rect 8008 -2139 8024 -2134
rect 8133 -2139 8135 -2099
rect 7813 -2323 8135 -2139
<< nsubdiff >>
rect 2991 -1619 3101 -1611
rect 2991 -1705 3003 -1619
rect 3089 -1705 3101 -1619
rect 2991 -1713 3101 -1705
<< nsubdiffcont >>
rect 3003 -1705 3089 -1619
<< locali >>
rect 275 625 1747 711
rect 275 371 361 625
rect 1661 585 1747 625
rect 1661 499 6685 585
rect 1735 465 2947 499
rect 3554 477 4643 499
rect -47 -85 39 64
rect 1103 -85 1189 45
rect -47 -101 1189 -85
rect -47 -135 409 -101
rect 443 -135 1189 -101
rect -47 -171 1189 -135
rect -148 -1294 -60 -1170
rect 2382 -1294 2470 -1170
rect -148 -1382 2470 -1294
rect 3020 -1354 3108 -1194
rect 5538 -1354 5626 -1212
rect 3020 -1442 5626 -1354
rect 6352 -1314 6440 -1166
rect 8878 -1314 8966 -1178
rect 6352 -1402 8966 -1314
rect 3003 -1616 3089 -1603
rect 3086 -1619 3089 -1616
rect 3086 -1707 3089 -1705
rect 3003 -4558 3089 -1707
rect 2556 -4580 4028 -4558
rect 2556 -4620 2580 -4580
rect 2620 -4620 4028 -4580
rect 2556 -4644 4028 -4620
<< viali >>
rect 555 415 589 449
rect 809 353 843 387
rect 409 229 443 263
rect 569 239 603 273
rect 2179 259 2213 293
rect 4119 265 4153 299
rect 6077 281 6111 315
rect 6320 214 6360 254
rect 409 -135 443 -101
rect 384 -1068 444 -1008
rect 1946 -1068 2006 -1008
rect 3444 -1110 3504 -1050
rect 5124 -1110 5184 -1050
rect 6755 -1079 6820 -1014
rect 8425 -1079 8491 -1013
rect 2995 -1619 3086 -1616
rect 2995 -1705 3003 -1619
rect 3003 -1705 3086 -1619
rect 2995 -1707 3086 -1705
rect 2580 -4620 2620 -4580
<< metal1 >>
rect 549 449 595 461
rect 549 415 555 449
rect 589 446 595 449
rect 589 418 840 446
rect 589 415 595 418
rect 549 403 595 415
rect 812 393 840 418
rect 803 387 849 393
rect 803 353 809 387
rect 843 353 849 387
rect 803 347 849 353
rect 6071 315 6117 321
rect 4107 299 4165 305
rect 2167 293 2225 299
rect 560 282 612 288
rect 397 263 455 269
rect 397 229 409 263
rect 443 229 455 263
rect 557 233 560 279
rect 397 223 455 229
rect 612 233 615 279
rect 2167 259 2179 293
rect 2213 259 2225 293
rect 4107 265 4119 299
rect 4153 298 4165 299
rect 4153 266 4232 298
rect 6071 281 6077 315
rect 6111 314 6117 315
rect 6111 282 6230 314
rect 6111 281 6117 282
rect 6071 275 6117 281
rect 4153 265 4165 266
rect 4107 259 4165 265
rect 2167 253 2225 259
rect 560 224 612 230
rect 410 -89 442 223
rect 403 -101 449 -89
rect 403 -135 409 -101
rect 443 -135 449 -101
rect 403 -147 449 -135
rect 2180 -294 2212 253
rect 1526 -326 2212 -294
rect 1526 -398 1558 -326
rect 4200 -390 4232 266
rect 4606 -390 4612 -380
rect 1516 -404 1568 -398
rect 4200 -422 4612 -390
rect 4606 -432 4612 -422
rect 4664 -432 4670 -380
rect 6198 -420 6230 282
rect 6308 208 6314 260
rect 6366 208 6372 260
rect 7960 -420 7966 -410
rect 6198 -452 7966 -420
rect 1516 -462 1568 -456
rect 7960 -462 7966 -452
rect 8018 -462 8024 -410
rect 378 -1008 450 -1002
rect 1940 -1008 2012 -996
rect -715 -1068 384 -1008
rect 444 -1068 1946 -1008
rect 2006 -1038 3504 -1008
rect 6749 -1013 6826 -1008
rect 8419 -1013 8497 -1007
rect 9578 -1013 9637 -1012
rect 6749 -1014 8425 -1013
rect 2006 -1050 3510 -1038
rect 5118 -1047 5190 -1044
rect 5922 -1047 5987 -1046
rect 6625 -1047 6755 -1014
rect 5118 -1050 6755 -1047
rect 2006 -1068 3444 -1050
rect -715 -1074 450 -1068
rect -715 -1076 448 -1074
rect -715 -4324 -647 -1076
rect 1940 -1080 2012 -1068
rect 824 -1956 884 -1950
rect 2688 -1956 2748 -1068
rect 3438 -1110 3444 -1068
rect 3504 -1110 5124 -1050
rect 5184 -1079 6755 -1050
rect 6820 -1079 8425 -1014
rect 8491 -1079 9258 -1013
rect 9482 -1072 10093 -1013
rect 9482 -1079 9541 -1072
rect 5184 -1110 6690 -1079
rect 6749 -1085 6826 -1079
rect 8419 -1085 8497 -1079
rect 3438 -1122 3510 -1110
rect 5118 -1112 6690 -1110
rect 5118 -1116 5190 -1112
rect 5922 -1289 5987 -1112
rect 5752 -1354 5987 -1289
rect 2983 -1616 3098 -1610
rect 2983 -1622 2995 -1616
rect 3086 -1622 3098 -1616
rect 2983 -1713 2989 -1622
rect 3092 -1713 3098 -1622
rect 2989 -1719 3092 -1713
rect 4618 -1871 4683 -1865
rect 5752 -1871 5817 -1354
rect 9578 -1738 9637 -1072
rect 4683 -1936 5817 -1871
rect 7943 -1797 9637 -1738
rect 4618 -1942 4683 -1936
rect 884 -2016 2748 -1956
rect 824 -2022 884 -2016
rect 7943 -2134 8002 -1797
rect 7943 -2199 8002 -2193
rect 9923 -4324 9978 -1072
rect -715 -4379 9978 -4324
rect -715 -4385 -647 -4379
rect 2574 -4574 2626 -4568
rect 2574 -4632 2626 -4626
<< via1 >>
rect 560 273 612 282
rect 560 239 569 273
rect 569 239 603 273
rect 603 239 612 273
rect 560 230 612 239
rect 1516 -456 1568 -404
rect 4612 -432 4664 -380
rect 6314 254 6366 260
rect 6314 214 6320 254
rect 6320 214 6360 254
rect 6360 214 6366 254
rect 6314 208 6366 214
rect 7966 -462 8018 -410
rect 2989 -1707 2995 -1622
rect 2995 -1707 3086 -1622
rect 3086 -1707 3092 -1622
rect 2989 -1713 3092 -1707
rect 4618 -1936 4683 -1871
rect 824 -2016 884 -1956
rect 7943 -2193 8002 -2134
rect 2574 -4580 2626 -4574
rect 2574 -4620 2580 -4580
rect 2580 -4620 2620 -4580
rect 2620 -4620 2626 -4580
rect 2574 -4626 2626 -4620
<< metal2 >>
rect 554 230 560 282
rect 612 230 618 282
rect 6314 260 6366 266
rect 570 -214 602 230
rect 6314 202 6366 208
rect 6324 -214 6356 202
rect 570 -246 6356 -214
rect 570 -518 602 -246
rect 4612 -376 4664 -374
rect 1510 -456 1512 -404
rect 1572 -456 1574 -404
rect 7966 -406 8018 -404
rect 4612 -438 4664 -436
rect 7966 -468 8018 -466
rect -344 -550 602 -518
rect -344 -4584 -312 -550
rect 2989 -1622 3092 -1613
rect 2983 -1713 2989 -1622
rect 3092 -1713 3098 -1622
rect 2989 -1722 3092 -1713
rect 4612 -1936 4618 -1871
rect 4683 -1936 4689 -1871
rect 818 -2016 824 -1956
rect 884 -2016 890 -1956
rect 7937 -2193 7943 -2134
rect 8003 -2193 8008 -2134
rect 2568 -4584 2574 -4574
rect -344 -4616 2574 -4584
rect 2568 -4626 2574 -4616
rect 2626 -4626 2632 -4574
<< via2 >>
rect 4608 -380 4668 -376
rect 1512 -404 1572 -400
rect 1512 -456 1516 -404
rect 1516 -456 1568 -404
rect 1568 -456 1572 -404
rect 4608 -432 4612 -380
rect 4612 -432 4664 -380
rect 4664 -432 4668 -380
rect 4608 -436 4668 -432
rect 7962 -410 8022 -406
rect 1512 -460 1572 -456
rect 7962 -462 7966 -410
rect 7966 -462 8018 -410
rect 8018 -462 8022 -410
rect 7962 -466 8022 -462
rect 9258 -1168 9482 -944
rect 2989 -1713 3092 -1622
rect 4618 -1936 4683 -1871
rect 824 -2016 884 -1956
rect 7943 -2134 8003 -2133
rect 7943 -2193 8002 -2134
rect 8002 -2193 8003 -2134
<< metal3 >>
rect 4612 -371 4812 -360
rect 4603 -376 4812 -371
rect 1507 -400 1577 -395
rect 1507 -404 1512 -400
rect 1456 -460 1512 -404
rect 1572 -404 1577 -400
rect 1572 -460 1656 -404
rect 4603 -436 4608 -376
rect 4668 -436 4812 -376
rect 7957 -406 8027 -401
rect 7957 -418 7962 -406
rect 4603 -441 4812 -436
rect 664 -1570 864 -1014
rect 1456 -1062 1656 -460
rect 4612 -1086 4812 -441
rect 7950 -466 7962 -418
rect 8022 -418 8027 -406
rect 8022 -466 8150 -418
rect 7950 -1058 8150 -466
rect 7164 -1570 7364 -1066
rect 664 -1770 2298 -1570
rect 2498 -1622 5932 -1570
rect 2498 -1713 2989 -1622
rect 3092 -1713 5932 -1622
rect 2498 -1770 5932 -1713
rect 6132 -1709 7364 -1570
rect 6132 -1770 7183 -1709
rect 7177 -1773 7183 -1770
rect 7417 -1773 7423 -1709
rect 819 -1956 889 -1951
rect 819 -1957 824 -1956
rect 884 -1957 889 -1956
rect 819 -2027 889 -2021
<< via3 >>
rect 2298 -1770 2498 -1570
rect 5932 -1770 6132 -1570
rect 7183 -1773 7417 -1709
rect 4613 -1871 4688 -1866
rect 4613 -1936 4618 -1871
rect 4618 -1936 4683 -1871
rect 4683 -1936 4688 -1871
rect 4613 -1941 4688 -1936
rect 819 -2016 824 -1957
rect 824 -2016 884 -1957
rect 884 -2016 889 -1957
rect 819 -2021 889 -2016
rect 7938 -2133 8008 -2128
rect 7938 -2193 7943 -2133
rect 7943 -2193 8003 -2133
rect 8003 -2193 8008 -2133
rect 7938 -2198 8008 -2193
<< via4 >>
rect 9252 -1174 9488 -938
rect 2238 -1570 2558 -1510
rect 2238 -1770 2298 -1570
rect 2298 -1770 2498 -1570
rect 2498 -1770 2558 -1570
rect 5872 -1570 6192 -1510
rect 694 -1957 1014 -1829
rect 2238 -1830 2558 -1770
rect 694 -2021 819 -1957
rect 819 -2021 889 -1957
rect 889 -2021 1014 -1957
rect 694 -2149 1014 -2021
rect 4491 -1866 4811 -1743
rect 5872 -1770 5932 -1570
rect 5932 -1770 6132 -1570
rect 6132 -1770 6192 -1570
rect 5872 -1830 6192 -1770
rect 7182 -1709 7418 -1538
rect 7182 -1773 7183 -1709
rect 7183 -1773 7417 -1709
rect 7417 -1773 7418 -1709
rect 7182 -1774 7418 -1773
rect 4491 -1941 4613 -1866
rect 4613 -1941 4688 -1866
rect 4688 -1941 4811 -1866
rect 4491 -2063 4811 -1941
rect 7813 -2128 8133 -2003
rect 7813 -2198 7938 -2128
rect 7938 -2198 8008 -2128
rect 8008 -2198 8133 -2128
rect 7813 -2323 8133 -2198
<< metal5 >>
rect 2214 -1510 2582 -1486
rect 670 -1829 1038 -1805
rect 670 -2149 694 -1829
rect 1014 -2149 1038 -1829
rect 2214 -1830 2238 -1510
rect 2558 -1830 2582 -1510
rect 5848 -1510 6216 -1486
rect 2214 -1854 2582 -1830
rect 4467 -1743 4835 -1719
rect 670 -2173 1038 -2149
rect 2238 -2156 2558 -1854
rect 4467 -2063 4491 -1743
rect 4811 -2063 4835 -1743
rect 5848 -1830 5872 -1510
rect 6192 -1830 6216 -1510
rect 7158 -1538 7442 -1514
rect 7158 -1774 7182 -1538
rect 7418 -1635 7442 -1538
rect 7418 -1677 9393 -1635
rect 7418 -1774 7442 -1677
rect 7158 -1798 7442 -1774
rect 5848 -1854 6216 -1830
rect 4467 -2087 4835 -2063
rect 694 -2314 1014 -2173
rect 4491 -2246 4811 -2087
rect 5872 -2138 6192 -1854
rect 7789 -2003 8157 -1979
rect 7789 -2323 7813 -2003
rect 8133 -2323 8157 -2003
rect 9351 -2060 9393 -1677
rect 7789 -2347 8157 -2323
use CNRATR_PCH_2C1F2  CNRATR_PCH_2C1F2_0 ~/aicex/ip/cnr_gr04_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 5502 0 1 60
box -184 -124 1336 613
use CNRATR_PCH_2C1F2  CNRATR_PCH_2C1F2_1
timestamp 1695852000
transform 1 0 -6 0 1 14
box -184 -124 1336 613
use CNRATR_PCH_2C1F2  CNRATR_PCH_2C1F2_2
timestamp 1695852000
transform 1 0 1764 0 1 26
box -184 -124 1336 613
use CNRATR_PCH_2C1F2  CNRATR_PCH_2C1F2_3
timestamp 1695852000
transform 1 0 3544 0 1 38
box -184 -124 1336 613
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_0
timestamp 1713472566
transform 1 0 8147 0 1 -3099
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_1
timestamp 1713472566
transform 1 0 1211 0 1 -3159
box -1349 -1081 1371 1081
use sky130_fd_pr__cap_mim_m3_2_KB5CJD  sky130_fd_pr__cap_mim_m3_2_KB5CJD_2
timestamp 1713472566
transform 1 0 4845 0 1 -3111
box -1349 -1081 1371 1081
use SUNTR_IVX1_CV  SUNTR_IVX1_CV_0 ~/aicex/ip/cnr_gr00_sky130nm/design/SUN_TR_SKY130NM
timestamp 1713466699
transform 1 0 6402 0 1 -1210
box -180 -132 2700 484
use SUNTR_IVX1_CV  SUNTR_IVX1_CV_1
timestamp 1713466699
transform 1 0 -92 0 1 -1214
box -180 -132 2700 484
use SUNTR_IVX1_CV  SUNTR_IVX1_CV_3
timestamp 1713466699
transform 1 0 3064 0 1 -1238
box -180 -132 2700 484
<< labels >>
flabel locali 275 625 1747 711 0 FreeSans 320 0 0 0 VDD_1V8
port 2 nsew
flabel locali 2556 -4644 4028 -4558 0 FreeSans 320 0 0 0 VSS
flabel metal1 9482 -1072 10093 -1013 0 FreeSans 320 0 0 0 OUT
port 4 nsew
<< end >>
